magic
tech sky130A
magscale 1 2
timestamp 1669602960
<< checkpaint >>
rect 512784 562457 515368 562502
rect 512721 559540 515401 562457
rect 512784 559460 515368 559540
<< error_p >>
rect 311757 484783 311793 484819
rect 283615 484699 283651 484735
rect 314281 482259 314317 482295
rect 281091 482175 281127 482211
rect 316805 479735 316841 479771
rect 278567 479651 278603 479687
rect 319329 477211 319365 477247
rect 276043 477127 276079 477163
rect 268722 472060 268758 472096
rect 263389 471887 263425 471923
rect 270286 470496 270322 470532
rect 265913 469363 265949 469399
rect 271850 468932 271886 468968
rect 268437 466839 268473 466875
rect 268437 464231 268473 464267
rect 271850 462114 271886 462150
rect 265913 461707 265949 461743
rect 270286 460550 270322 460586
rect 263389 459183 263425 459219
rect 268722 458986 268758 459022
rect 276063 453907 276099 453943
rect 319332 453823 319368 453859
rect 278587 451383 278623 451419
rect 316808 451299 316844 451335
rect 281111 448859 281147 448895
rect 314284 448775 314320 448811
rect 283635 446335 283671 446371
rect 311760 446251 311796 446287
rect 452088 332526 452090 373009
rect 454892 366099 454893 373009
rect 455012 366183 455013 373009
rect 452288 363324 452289 366099
rect 454893 362417 454894 365891
rect 455013 362537 455014 365891
rect 452090 320998 452091 331259
rect 452289 317354 452291 362417
<< error_s >>
rect 152640 437073 152653 437237
rect 163097 437229 163105 437237
rect 163105 437209 163116 437229
rect 152334 436926 152481 436929
rect 152318 436777 152334 436926
rect 163441 436873 163461 436875
rect 163461 436865 163469 436873
rect 163469 436845 163478 436865
rect 152014 436606 152185 436609
rect 151998 436513 152014 436606
rect 163777 436552 163782 436555
rect 163782 436529 163798 436552
rect 151694 436286 151914 436289
rect 151678 436053 151694 436286
rect 163882 436232 164102 436235
rect 164102 435999 164118 436232
rect 151371 435963 151591 435966
rect 151355 435939 151371 435963
rect 468118 428041 468688 428060
rect 481206 428041 481776 428060
rect 411902 428021 412472 428040
rect 424990 428021 425560 428040
rect 425892 428021 426462 428040
rect 438980 428021 439550 428040
rect 439882 428021 440452 428040
rect 452970 428021 453540 428040
rect 456242 428021 456812 428040
rect 411902 427627 412489 428021
rect 424990 427627 425577 428021
rect 425892 427627 426479 428021
rect 438980 427627 439567 428021
rect 439882 427627 440469 428021
rect 452970 427627 453557 428021
rect 456242 427627 456829 428021
rect 468118 427647 468705 428041
rect 481206 427647 481793 428041
rect 468118 427628 468688 427647
rect 481206 427628 481776 427647
rect 411902 427608 412472 427627
rect 424990 427608 425560 427627
rect 425892 427608 426462 427627
rect 438980 427608 439550 427627
rect 439882 427608 440452 427627
rect 452970 427608 453540 427627
rect 456242 427608 456812 427627
rect 468118 427276 468688 427296
rect 469754 427276 470324 427296
rect 471390 427276 471960 427296
rect 473026 427276 473596 427296
rect 474662 427276 475232 427296
rect 476298 427276 476868 427296
rect 416810 427256 417380 427276
rect 418446 427256 419016 427276
rect 420082 427256 420652 427276
rect 421718 427256 422288 427276
rect 423354 427256 423924 427276
rect 424990 427256 425560 427276
rect 430800 427256 431370 427276
rect 432436 427256 433006 427276
rect 434072 427256 434642 427276
rect 435708 427256 436278 427276
rect 437344 427256 437914 427276
rect 438980 427256 439550 427276
rect 444790 427256 445360 427276
rect 446426 427256 446996 427276
rect 448062 427256 448632 427276
rect 449698 427256 450268 427276
rect 451334 427256 451904 427276
rect 452970 427256 453540 427276
rect 454606 427256 455176 427276
rect 456242 427256 456812 427276
rect 416810 426862 417397 427256
rect 418446 426862 419033 427256
rect 420082 426862 420669 427256
rect 421718 426862 422305 427256
rect 423354 426862 423941 427256
rect 424990 426862 425577 427256
rect 430800 426862 431387 427256
rect 432436 426862 433023 427256
rect 434072 426862 434659 427256
rect 435708 426862 436295 427256
rect 437344 426862 437931 427256
rect 438980 426862 439567 427256
rect 444790 426862 445377 427256
rect 446426 426862 447013 427256
rect 448062 426862 448649 427256
rect 449698 426862 450285 427256
rect 451334 426862 451921 427256
rect 452970 426862 453557 427256
rect 454606 426862 455193 427256
rect 456242 426862 456829 427256
rect 468118 426882 468705 427276
rect 469754 426882 470341 427276
rect 471390 426882 471977 427276
rect 473026 426882 473613 427276
rect 474662 426882 475249 427276
rect 476298 426882 476885 427276
rect 468118 426864 468688 426882
rect 469754 426864 470324 426882
rect 471390 426864 471960 426882
rect 473026 426864 473596 426882
rect 474662 426864 475232 426882
rect 476298 426864 476868 426882
rect 416810 426844 417380 426862
rect 418446 426844 419016 426862
rect 420082 426844 420652 426862
rect 421718 426844 422288 426862
rect 423354 426844 423924 426862
rect 424990 426844 425560 426862
rect 430800 426844 431370 426862
rect 432436 426844 433006 426862
rect 434072 426844 434642 426862
rect 435708 426844 436278 426862
rect 437344 426844 437914 426862
rect 438980 426844 439550 426862
rect 444790 426844 445360 426862
rect 446426 426844 446996 426862
rect 448062 426844 448632 426862
rect 449698 426844 450268 426862
rect 451334 426844 451904 426862
rect 452970 426844 453540 426862
rect 454606 426844 455176 426862
rect 456242 426844 456812 426862
rect 164371 423479 164387 423503
rect 164151 423476 164371 423479
rect 151624 423210 151640 423443
rect 151640 423207 151860 423210
rect 164048 423156 164064 423243
rect 163853 423153 164048 423156
rect 151944 422890 151960 422983
rect 151960 422887 152180 422890
rect 163741 422849 163744 422877
rect 163713 422833 163741 422849
rect 152264 422570 152280 422665
rect 152280 422567 152399 422570
rect 163408 422516 163424 422541
rect 163405 422513 163408 422516
rect 152626 422208 152642 422441
rect 152642 422205 152653 422208
rect 163097 422205 163102 422233
rect 152640 299523 152653 299687
rect 163097 299679 163105 299687
rect 163105 299659 163116 299679
rect 152334 299376 152481 299379
rect 152318 299227 152334 299376
rect 163441 299323 163461 299325
rect 163461 299315 163469 299323
rect 163469 299295 163478 299315
rect 152014 299056 152185 299059
rect 151998 298963 152014 299056
rect 163777 299002 163782 299005
rect 163782 298979 163798 299002
rect 151694 298736 151914 298739
rect 151678 298503 151694 298736
rect 163882 298682 164102 298685
rect 164102 298449 164118 298682
rect 151371 298413 151591 298416
rect 151355 298389 151371 298413
rect 164371 285929 164387 285953
rect 164151 285926 164371 285929
rect 151624 285660 151640 285893
rect 151640 285657 151860 285660
rect 164048 285606 164064 285693
rect 163853 285603 164048 285606
rect 151944 285340 151960 285433
rect 151960 285337 152180 285340
rect 163741 285299 163744 285327
rect 163713 285283 163741 285299
rect 152264 285020 152280 285115
rect 152280 285017 152399 285020
rect 163408 284966 163424 284991
rect 163405 284963 163408 284966
rect 152626 284658 152642 284891
rect 152642 284655 152653 284658
rect 163097 284655 163102 284683
<< dnwell >>
rect 10605 686997 12505 688897
rect 10605 683750 12505 685650
rect 509057 555465 510957 557365
rect 514903 555465 516803 557365
rect 151045 420664 164835 447064
rect 151045 283114 164835 309514
<< nwell >>
rect 508977 557159 511037 557445
rect 508977 555671 509263 557159
rect 510751 555671 511037 557159
rect 508977 555385 511037 555671
rect 514823 557159 516883 557445
rect 514823 555671 515109 557159
rect 516597 555671 516883 557159
rect 514823 555385 516883 555671
<< pwell >>
rect 509467 557599 510523 558655
rect 515313 557599 516369 558655
rect 509467 555899 510523 556955
rect 515313 555899 516369 556955
<< psubdiff >>
rect 509493 558595 509604 558629
rect 509638 558595 509672 558629
rect 509706 558595 509740 558629
rect 509774 558595 509808 558629
rect 509842 558595 509876 558629
rect 509910 558595 509944 558629
rect 509978 558595 510012 558629
rect 510046 558595 510080 558629
rect 510114 558595 510148 558629
rect 510182 558595 510216 558629
rect 510250 558595 510284 558629
rect 510318 558595 510352 558629
rect 510386 558595 510497 558629
rect 509493 558518 509527 558595
rect 509493 558450 509527 558484
rect 509493 558382 509527 558416
rect 509493 558314 509527 558348
rect 509493 558246 509527 558280
rect 509493 558178 509527 558212
rect 509493 558110 509527 558144
rect 509493 558042 509527 558076
rect 509493 557974 509527 558008
rect 509493 557906 509527 557940
rect 509493 557838 509527 557872
rect 509493 557770 509527 557804
rect 509493 557659 509527 557736
rect 510463 558518 510497 558595
rect 510463 558450 510497 558484
rect 510463 558382 510497 558416
rect 510463 558314 510497 558348
rect 510463 558246 510497 558280
rect 510463 558178 510497 558212
rect 510463 558110 510497 558144
rect 510463 558042 510497 558076
rect 510463 557974 510497 558008
rect 510463 557906 510497 557940
rect 510463 557838 510497 557872
rect 510463 557770 510497 557804
rect 510463 557659 510497 557736
rect 509493 557625 509604 557659
rect 509638 557625 509672 557659
rect 509706 557625 509740 557659
rect 509774 557625 509808 557659
rect 509842 557625 509876 557659
rect 509910 557625 509944 557659
rect 509978 557625 510012 557659
rect 510046 557625 510080 557659
rect 510114 557625 510148 557659
rect 510182 557625 510216 557659
rect 510250 557625 510284 557659
rect 510318 557625 510352 557659
rect 510386 557625 510497 557659
rect 515339 558595 515450 558629
rect 515484 558595 515518 558629
rect 515552 558595 515586 558629
rect 515620 558595 515654 558629
rect 515688 558595 515722 558629
rect 515756 558595 515790 558629
rect 515824 558595 515858 558629
rect 515892 558595 515926 558629
rect 515960 558595 515994 558629
rect 516028 558595 516062 558629
rect 516096 558595 516130 558629
rect 516164 558595 516198 558629
rect 516232 558595 516343 558629
rect 515339 558518 515373 558595
rect 515339 558450 515373 558484
rect 515339 558382 515373 558416
rect 515339 558314 515373 558348
rect 515339 558246 515373 558280
rect 515339 558178 515373 558212
rect 515339 558110 515373 558144
rect 515339 558042 515373 558076
rect 515339 557974 515373 558008
rect 515339 557906 515373 557940
rect 515339 557838 515373 557872
rect 515339 557770 515373 557804
rect 515339 557659 515373 557736
rect 516309 558518 516343 558595
rect 516309 558450 516343 558484
rect 516309 558382 516343 558416
rect 516309 558314 516343 558348
rect 516309 558246 516343 558280
rect 516309 558178 516343 558212
rect 516309 558110 516343 558144
rect 516309 558042 516343 558076
rect 516309 557974 516343 558008
rect 516309 557906 516343 557940
rect 516309 557838 516343 557872
rect 516309 557770 516343 557804
rect 516309 557659 516343 557736
rect 515339 557625 515450 557659
rect 515484 557625 515518 557659
rect 515552 557625 515586 557659
rect 515620 557625 515654 557659
rect 515688 557625 515722 557659
rect 515756 557625 515790 557659
rect 515824 557625 515858 557659
rect 515892 557625 515926 557659
rect 515960 557625 515994 557659
rect 516028 557625 516062 557659
rect 516096 557625 516130 557659
rect 516164 557625 516198 557659
rect 516232 557625 516343 557659
rect 509493 556895 509604 556929
rect 509638 556895 509672 556929
rect 509706 556895 509740 556929
rect 509774 556895 509808 556929
rect 509842 556895 509876 556929
rect 509910 556895 509944 556929
rect 509978 556895 510012 556929
rect 510046 556895 510080 556929
rect 510114 556895 510148 556929
rect 510182 556895 510216 556929
rect 510250 556895 510284 556929
rect 510318 556895 510352 556929
rect 510386 556895 510497 556929
rect 509493 556818 509527 556895
rect 509493 556750 509527 556784
rect 509493 556682 509527 556716
rect 509493 556614 509527 556648
rect 509493 556546 509527 556580
rect 509493 556478 509527 556512
rect 509493 556410 509527 556444
rect 509493 556342 509527 556376
rect 509493 556274 509527 556308
rect 509493 556206 509527 556240
rect 509493 556138 509527 556172
rect 509493 556070 509527 556104
rect 509493 555959 509527 556036
rect 510463 556818 510497 556895
rect 510463 556750 510497 556784
rect 510463 556682 510497 556716
rect 510463 556614 510497 556648
rect 510463 556546 510497 556580
rect 510463 556478 510497 556512
rect 510463 556410 510497 556444
rect 510463 556342 510497 556376
rect 510463 556274 510497 556308
rect 510463 556206 510497 556240
rect 510463 556138 510497 556172
rect 510463 556070 510497 556104
rect 510463 555959 510497 556036
rect 509493 555925 509604 555959
rect 509638 555925 509672 555959
rect 509706 555925 509740 555959
rect 509774 555925 509808 555959
rect 509842 555925 509876 555959
rect 509910 555925 509944 555959
rect 509978 555925 510012 555959
rect 510046 555925 510080 555959
rect 510114 555925 510148 555959
rect 510182 555925 510216 555959
rect 510250 555925 510284 555959
rect 510318 555925 510352 555959
rect 510386 555925 510497 555959
rect 515339 556895 515450 556929
rect 515484 556895 515518 556929
rect 515552 556895 515586 556929
rect 515620 556895 515654 556929
rect 515688 556895 515722 556929
rect 515756 556895 515790 556929
rect 515824 556895 515858 556929
rect 515892 556895 515926 556929
rect 515960 556895 515994 556929
rect 516028 556895 516062 556929
rect 516096 556895 516130 556929
rect 516164 556895 516198 556929
rect 516232 556895 516343 556929
rect 515339 556818 515373 556895
rect 515339 556750 515373 556784
rect 515339 556682 515373 556716
rect 515339 556614 515373 556648
rect 515339 556546 515373 556580
rect 515339 556478 515373 556512
rect 515339 556410 515373 556444
rect 515339 556342 515373 556376
rect 515339 556274 515373 556308
rect 515339 556206 515373 556240
rect 515339 556138 515373 556172
rect 515339 556070 515373 556104
rect 515339 555959 515373 556036
rect 516309 556818 516343 556895
rect 516309 556750 516343 556784
rect 516309 556682 516343 556716
rect 516309 556614 516343 556648
rect 516309 556546 516343 556580
rect 516309 556478 516343 556512
rect 516309 556410 516343 556444
rect 516309 556342 516343 556376
rect 516309 556274 516343 556308
rect 516309 556206 516343 556240
rect 516309 556138 516343 556172
rect 516309 556070 516343 556104
rect 516309 555959 516343 556036
rect 515339 555925 515450 555959
rect 515484 555925 515518 555959
rect 515552 555925 515586 555959
rect 515620 555925 515654 555959
rect 515688 555925 515722 555959
rect 515756 555925 515790 555959
rect 515824 555925 515858 555959
rect 515892 555925 515926 555959
rect 515960 555925 515994 555959
rect 516028 555925 516062 555959
rect 516096 555925 516130 555959
rect 516164 555925 516198 555959
rect 516232 555925 516343 555959
<< nsubdiff >>
rect 509014 557388 511000 557408
rect 509014 557354 509106 557388
rect 509140 557354 509174 557388
rect 509208 557354 509242 557388
rect 509276 557354 509310 557388
rect 509344 557354 509378 557388
rect 509412 557354 509446 557388
rect 509480 557354 509514 557388
rect 509548 557354 509582 557388
rect 509616 557354 509650 557388
rect 509684 557354 509718 557388
rect 509752 557354 509786 557388
rect 509820 557354 509854 557388
rect 509888 557354 509922 557388
rect 509956 557354 509990 557388
rect 510024 557354 510058 557388
rect 510092 557354 510126 557388
rect 510160 557354 510194 557388
rect 510228 557354 510262 557388
rect 510296 557354 510330 557388
rect 510364 557354 510398 557388
rect 510432 557354 510466 557388
rect 510500 557354 510534 557388
rect 510568 557354 510602 557388
rect 510636 557354 510670 557388
rect 510704 557354 510738 557388
rect 510772 557354 510806 557388
rect 510840 557354 510874 557388
rect 510908 557354 511000 557388
rect 509014 557334 511000 557354
rect 509014 557316 509088 557334
rect 509014 557282 509034 557316
rect 509068 557282 509088 557316
rect 509014 557248 509088 557282
rect 509014 557214 509034 557248
rect 509068 557214 509088 557248
rect 509014 557180 509088 557214
rect 509014 557146 509034 557180
rect 509068 557146 509088 557180
rect 509014 557112 509088 557146
rect 509014 557078 509034 557112
rect 509068 557078 509088 557112
rect 509014 557044 509088 557078
rect 509014 557010 509034 557044
rect 509068 557010 509088 557044
rect 509014 556976 509088 557010
rect 509014 556942 509034 556976
rect 509068 556942 509088 556976
rect 509014 556908 509088 556942
rect 510926 557316 511000 557334
rect 510926 557282 510946 557316
rect 510980 557282 511000 557316
rect 510926 557248 511000 557282
rect 510926 557214 510946 557248
rect 510980 557214 511000 557248
rect 510926 557180 511000 557214
rect 510926 557146 510946 557180
rect 510980 557146 511000 557180
rect 510926 557112 511000 557146
rect 510926 557078 510946 557112
rect 510980 557078 511000 557112
rect 510926 557044 511000 557078
rect 510926 557010 510946 557044
rect 510980 557010 511000 557044
rect 510926 556976 511000 557010
rect 510926 556942 510946 556976
rect 510980 556942 511000 556976
rect 509014 556874 509034 556908
rect 509068 556874 509088 556908
rect 509014 556840 509088 556874
rect 509014 556806 509034 556840
rect 509068 556806 509088 556840
rect 509014 556772 509088 556806
rect 509014 556738 509034 556772
rect 509068 556738 509088 556772
rect 509014 556704 509088 556738
rect 509014 556670 509034 556704
rect 509068 556670 509088 556704
rect 509014 556636 509088 556670
rect 509014 556602 509034 556636
rect 509068 556602 509088 556636
rect 509014 556568 509088 556602
rect 509014 556534 509034 556568
rect 509068 556534 509088 556568
rect 509014 556500 509088 556534
rect 509014 556466 509034 556500
rect 509068 556466 509088 556500
rect 509014 556432 509088 556466
rect 509014 556398 509034 556432
rect 509068 556398 509088 556432
rect 509014 556364 509088 556398
rect 509014 556330 509034 556364
rect 509068 556330 509088 556364
rect 509014 556296 509088 556330
rect 509014 556262 509034 556296
rect 509068 556262 509088 556296
rect 509014 556228 509088 556262
rect 509014 556194 509034 556228
rect 509068 556194 509088 556228
rect 509014 556160 509088 556194
rect 509014 556126 509034 556160
rect 509068 556126 509088 556160
rect 509014 556092 509088 556126
rect 509014 556058 509034 556092
rect 509068 556058 509088 556092
rect 509014 556024 509088 556058
rect 509014 555990 509034 556024
rect 509068 555990 509088 556024
rect 509014 555956 509088 555990
rect 509014 555922 509034 555956
rect 509068 555922 509088 555956
rect 510926 556908 511000 556942
rect 510926 556874 510946 556908
rect 510980 556874 511000 556908
rect 510926 556840 511000 556874
rect 510926 556806 510946 556840
rect 510980 556806 511000 556840
rect 510926 556772 511000 556806
rect 510926 556738 510946 556772
rect 510980 556738 511000 556772
rect 510926 556704 511000 556738
rect 510926 556670 510946 556704
rect 510980 556670 511000 556704
rect 510926 556636 511000 556670
rect 510926 556602 510946 556636
rect 510980 556602 511000 556636
rect 510926 556568 511000 556602
rect 510926 556534 510946 556568
rect 510980 556534 511000 556568
rect 510926 556500 511000 556534
rect 510926 556466 510946 556500
rect 510980 556466 511000 556500
rect 510926 556432 511000 556466
rect 510926 556398 510946 556432
rect 510980 556398 511000 556432
rect 510926 556364 511000 556398
rect 510926 556330 510946 556364
rect 510980 556330 511000 556364
rect 510926 556296 511000 556330
rect 510926 556262 510946 556296
rect 510980 556262 511000 556296
rect 510926 556228 511000 556262
rect 510926 556194 510946 556228
rect 510980 556194 511000 556228
rect 510926 556160 511000 556194
rect 510926 556126 510946 556160
rect 510980 556126 511000 556160
rect 510926 556092 511000 556126
rect 510926 556058 510946 556092
rect 510980 556058 511000 556092
rect 510926 556024 511000 556058
rect 510926 555990 510946 556024
rect 510980 555990 511000 556024
rect 510926 555956 511000 555990
rect 509014 555888 509088 555922
rect 509014 555854 509034 555888
rect 509068 555854 509088 555888
rect 509014 555820 509088 555854
rect 509014 555786 509034 555820
rect 509068 555786 509088 555820
rect 509014 555752 509088 555786
rect 509014 555718 509034 555752
rect 509068 555718 509088 555752
rect 509014 555684 509088 555718
rect 509014 555650 509034 555684
rect 509068 555650 509088 555684
rect 509014 555616 509088 555650
rect 509014 555582 509034 555616
rect 509068 555582 509088 555616
rect 509014 555548 509088 555582
rect 509014 555514 509034 555548
rect 509068 555514 509088 555548
rect 509014 555496 509088 555514
rect 510926 555922 510946 555956
rect 510980 555922 511000 555956
rect 510926 555888 511000 555922
rect 510926 555854 510946 555888
rect 510980 555854 511000 555888
rect 510926 555820 511000 555854
rect 510926 555786 510946 555820
rect 510980 555786 511000 555820
rect 510926 555752 511000 555786
rect 510926 555718 510946 555752
rect 510980 555718 511000 555752
rect 510926 555684 511000 555718
rect 510926 555650 510946 555684
rect 510980 555650 511000 555684
rect 510926 555616 511000 555650
rect 510926 555582 510946 555616
rect 510980 555582 511000 555616
rect 510926 555548 511000 555582
rect 510926 555514 510946 555548
rect 510980 555514 511000 555548
rect 510926 555496 511000 555514
rect 509014 555476 511000 555496
rect 509014 555442 509106 555476
rect 509140 555442 509174 555476
rect 509208 555442 509242 555476
rect 509276 555442 509310 555476
rect 509344 555442 509378 555476
rect 509412 555442 509446 555476
rect 509480 555442 509514 555476
rect 509548 555442 509582 555476
rect 509616 555442 509650 555476
rect 509684 555442 509718 555476
rect 509752 555442 509786 555476
rect 509820 555442 509854 555476
rect 509888 555442 509922 555476
rect 509956 555442 509990 555476
rect 510024 555442 510058 555476
rect 510092 555442 510126 555476
rect 510160 555442 510194 555476
rect 510228 555442 510262 555476
rect 510296 555442 510330 555476
rect 510364 555442 510398 555476
rect 510432 555442 510466 555476
rect 510500 555442 510534 555476
rect 510568 555442 510602 555476
rect 510636 555442 510670 555476
rect 510704 555442 510738 555476
rect 510772 555442 510806 555476
rect 510840 555442 510874 555476
rect 510908 555442 511000 555476
rect 509014 555422 511000 555442
rect 514860 557388 516846 557408
rect 514860 557354 514952 557388
rect 514986 557354 515020 557388
rect 515054 557354 515088 557388
rect 515122 557354 515156 557388
rect 515190 557354 515224 557388
rect 515258 557354 515292 557388
rect 515326 557354 515360 557388
rect 515394 557354 515428 557388
rect 515462 557354 515496 557388
rect 515530 557354 515564 557388
rect 515598 557354 515632 557388
rect 515666 557354 515700 557388
rect 515734 557354 515768 557388
rect 515802 557354 515836 557388
rect 515870 557354 515904 557388
rect 515938 557354 515972 557388
rect 516006 557354 516040 557388
rect 516074 557354 516108 557388
rect 516142 557354 516176 557388
rect 516210 557354 516244 557388
rect 516278 557354 516312 557388
rect 516346 557354 516380 557388
rect 516414 557354 516448 557388
rect 516482 557354 516516 557388
rect 516550 557354 516584 557388
rect 516618 557354 516652 557388
rect 516686 557354 516720 557388
rect 516754 557354 516846 557388
rect 514860 557334 516846 557354
rect 514860 557316 514934 557334
rect 514860 557282 514880 557316
rect 514914 557282 514934 557316
rect 514860 557248 514934 557282
rect 514860 557214 514880 557248
rect 514914 557214 514934 557248
rect 514860 557180 514934 557214
rect 514860 557146 514880 557180
rect 514914 557146 514934 557180
rect 514860 557112 514934 557146
rect 514860 557078 514880 557112
rect 514914 557078 514934 557112
rect 514860 557044 514934 557078
rect 514860 557010 514880 557044
rect 514914 557010 514934 557044
rect 514860 556976 514934 557010
rect 514860 556942 514880 556976
rect 514914 556942 514934 556976
rect 514860 556908 514934 556942
rect 516772 557316 516846 557334
rect 516772 557282 516792 557316
rect 516826 557282 516846 557316
rect 516772 557248 516846 557282
rect 516772 557214 516792 557248
rect 516826 557214 516846 557248
rect 516772 557180 516846 557214
rect 516772 557146 516792 557180
rect 516826 557146 516846 557180
rect 516772 557112 516846 557146
rect 516772 557078 516792 557112
rect 516826 557078 516846 557112
rect 516772 557044 516846 557078
rect 516772 557010 516792 557044
rect 516826 557010 516846 557044
rect 516772 556976 516846 557010
rect 516772 556942 516792 556976
rect 516826 556942 516846 556976
rect 514860 556874 514880 556908
rect 514914 556874 514934 556908
rect 514860 556840 514934 556874
rect 514860 556806 514880 556840
rect 514914 556806 514934 556840
rect 514860 556772 514934 556806
rect 514860 556738 514880 556772
rect 514914 556738 514934 556772
rect 514860 556704 514934 556738
rect 514860 556670 514880 556704
rect 514914 556670 514934 556704
rect 514860 556636 514934 556670
rect 514860 556602 514880 556636
rect 514914 556602 514934 556636
rect 514860 556568 514934 556602
rect 514860 556534 514880 556568
rect 514914 556534 514934 556568
rect 514860 556500 514934 556534
rect 514860 556466 514880 556500
rect 514914 556466 514934 556500
rect 514860 556432 514934 556466
rect 514860 556398 514880 556432
rect 514914 556398 514934 556432
rect 514860 556364 514934 556398
rect 514860 556330 514880 556364
rect 514914 556330 514934 556364
rect 514860 556296 514934 556330
rect 514860 556262 514880 556296
rect 514914 556262 514934 556296
rect 514860 556228 514934 556262
rect 514860 556194 514880 556228
rect 514914 556194 514934 556228
rect 514860 556160 514934 556194
rect 514860 556126 514880 556160
rect 514914 556126 514934 556160
rect 514860 556092 514934 556126
rect 514860 556058 514880 556092
rect 514914 556058 514934 556092
rect 514860 556024 514934 556058
rect 514860 555990 514880 556024
rect 514914 555990 514934 556024
rect 514860 555956 514934 555990
rect 514860 555922 514880 555956
rect 514914 555922 514934 555956
rect 516772 556908 516846 556942
rect 516772 556874 516792 556908
rect 516826 556874 516846 556908
rect 516772 556840 516846 556874
rect 516772 556806 516792 556840
rect 516826 556806 516846 556840
rect 516772 556772 516846 556806
rect 516772 556738 516792 556772
rect 516826 556738 516846 556772
rect 516772 556704 516846 556738
rect 516772 556670 516792 556704
rect 516826 556670 516846 556704
rect 516772 556636 516846 556670
rect 516772 556602 516792 556636
rect 516826 556602 516846 556636
rect 516772 556568 516846 556602
rect 516772 556534 516792 556568
rect 516826 556534 516846 556568
rect 516772 556500 516846 556534
rect 516772 556466 516792 556500
rect 516826 556466 516846 556500
rect 516772 556432 516846 556466
rect 516772 556398 516792 556432
rect 516826 556398 516846 556432
rect 516772 556364 516846 556398
rect 516772 556330 516792 556364
rect 516826 556330 516846 556364
rect 516772 556296 516846 556330
rect 516772 556262 516792 556296
rect 516826 556262 516846 556296
rect 516772 556228 516846 556262
rect 516772 556194 516792 556228
rect 516826 556194 516846 556228
rect 516772 556160 516846 556194
rect 516772 556126 516792 556160
rect 516826 556126 516846 556160
rect 516772 556092 516846 556126
rect 516772 556058 516792 556092
rect 516826 556058 516846 556092
rect 516772 556024 516846 556058
rect 516772 555990 516792 556024
rect 516826 555990 516846 556024
rect 516772 555956 516846 555990
rect 514860 555888 514934 555922
rect 514860 555854 514880 555888
rect 514914 555854 514934 555888
rect 514860 555820 514934 555854
rect 514860 555786 514880 555820
rect 514914 555786 514934 555820
rect 514860 555752 514934 555786
rect 514860 555718 514880 555752
rect 514914 555718 514934 555752
rect 514860 555684 514934 555718
rect 514860 555650 514880 555684
rect 514914 555650 514934 555684
rect 514860 555616 514934 555650
rect 514860 555582 514880 555616
rect 514914 555582 514934 555616
rect 514860 555548 514934 555582
rect 514860 555514 514880 555548
rect 514914 555514 514934 555548
rect 514860 555496 514934 555514
rect 516772 555922 516792 555956
rect 516826 555922 516846 555956
rect 516772 555888 516846 555922
rect 516772 555854 516792 555888
rect 516826 555854 516846 555888
rect 516772 555820 516846 555854
rect 516772 555786 516792 555820
rect 516826 555786 516846 555820
rect 516772 555752 516846 555786
rect 516772 555718 516792 555752
rect 516826 555718 516846 555752
rect 516772 555684 516846 555718
rect 516772 555650 516792 555684
rect 516826 555650 516846 555684
rect 516772 555616 516846 555650
rect 516772 555582 516792 555616
rect 516826 555582 516846 555616
rect 516772 555548 516846 555582
rect 516772 555514 516792 555548
rect 516826 555514 516846 555548
rect 516772 555496 516846 555514
rect 514860 555476 516846 555496
rect 514860 555442 514952 555476
rect 514986 555442 515020 555476
rect 515054 555442 515088 555476
rect 515122 555442 515156 555476
rect 515190 555442 515224 555476
rect 515258 555442 515292 555476
rect 515326 555442 515360 555476
rect 515394 555442 515428 555476
rect 515462 555442 515496 555476
rect 515530 555442 515564 555476
rect 515598 555442 515632 555476
rect 515666 555442 515700 555476
rect 515734 555442 515768 555476
rect 515802 555442 515836 555476
rect 515870 555442 515904 555476
rect 515938 555442 515972 555476
rect 516006 555442 516040 555476
rect 516074 555442 516108 555476
rect 516142 555442 516176 555476
rect 516210 555442 516244 555476
rect 516278 555442 516312 555476
rect 516346 555442 516380 555476
rect 516414 555442 516448 555476
rect 516482 555442 516516 555476
rect 516550 555442 516584 555476
rect 516618 555442 516652 555476
rect 516686 555442 516720 555476
rect 516754 555442 516846 555476
rect 514860 555422 516846 555442
<< psubdiffcont >>
rect 509604 558595 509638 558629
rect 509672 558595 509706 558629
rect 509740 558595 509774 558629
rect 509808 558595 509842 558629
rect 509876 558595 509910 558629
rect 509944 558595 509978 558629
rect 510012 558595 510046 558629
rect 510080 558595 510114 558629
rect 510148 558595 510182 558629
rect 510216 558595 510250 558629
rect 510284 558595 510318 558629
rect 510352 558595 510386 558629
rect 509493 558484 509527 558518
rect 509493 558416 509527 558450
rect 509493 558348 509527 558382
rect 509493 558280 509527 558314
rect 509493 558212 509527 558246
rect 509493 558144 509527 558178
rect 509493 558076 509527 558110
rect 509493 558008 509527 558042
rect 509493 557940 509527 557974
rect 509493 557872 509527 557906
rect 509493 557804 509527 557838
rect 509493 557736 509527 557770
rect 510463 558484 510497 558518
rect 510463 558416 510497 558450
rect 510463 558348 510497 558382
rect 510463 558280 510497 558314
rect 510463 558212 510497 558246
rect 510463 558144 510497 558178
rect 510463 558076 510497 558110
rect 510463 558008 510497 558042
rect 510463 557940 510497 557974
rect 510463 557872 510497 557906
rect 510463 557804 510497 557838
rect 510463 557736 510497 557770
rect 509604 557625 509638 557659
rect 509672 557625 509706 557659
rect 509740 557625 509774 557659
rect 509808 557625 509842 557659
rect 509876 557625 509910 557659
rect 509944 557625 509978 557659
rect 510012 557625 510046 557659
rect 510080 557625 510114 557659
rect 510148 557625 510182 557659
rect 510216 557625 510250 557659
rect 510284 557625 510318 557659
rect 510352 557625 510386 557659
rect 515450 558595 515484 558629
rect 515518 558595 515552 558629
rect 515586 558595 515620 558629
rect 515654 558595 515688 558629
rect 515722 558595 515756 558629
rect 515790 558595 515824 558629
rect 515858 558595 515892 558629
rect 515926 558595 515960 558629
rect 515994 558595 516028 558629
rect 516062 558595 516096 558629
rect 516130 558595 516164 558629
rect 516198 558595 516232 558629
rect 515339 558484 515373 558518
rect 515339 558416 515373 558450
rect 515339 558348 515373 558382
rect 515339 558280 515373 558314
rect 515339 558212 515373 558246
rect 515339 558144 515373 558178
rect 515339 558076 515373 558110
rect 515339 558008 515373 558042
rect 515339 557940 515373 557974
rect 515339 557872 515373 557906
rect 515339 557804 515373 557838
rect 515339 557736 515373 557770
rect 516309 558484 516343 558518
rect 516309 558416 516343 558450
rect 516309 558348 516343 558382
rect 516309 558280 516343 558314
rect 516309 558212 516343 558246
rect 516309 558144 516343 558178
rect 516309 558076 516343 558110
rect 516309 558008 516343 558042
rect 516309 557940 516343 557974
rect 516309 557872 516343 557906
rect 516309 557804 516343 557838
rect 516309 557736 516343 557770
rect 515450 557625 515484 557659
rect 515518 557625 515552 557659
rect 515586 557625 515620 557659
rect 515654 557625 515688 557659
rect 515722 557625 515756 557659
rect 515790 557625 515824 557659
rect 515858 557625 515892 557659
rect 515926 557625 515960 557659
rect 515994 557625 516028 557659
rect 516062 557625 516096 557659
rect 516130 557625 516164 557659
rect 516198 557625 516232 557659
rect 509604 556895 509638 556929
rect 509672 556895 509706 556929
rect 509740 556895 509774 556929
rect 509808 556895 509842 556929
rect 509876 556895 509910 556929
rect 509944 556895 509978 556929
rect 510012 556895 510046 556929
rect 510080 556895 510114 556929
rect 510148 556895 510182 556929
rect 510216 556895 510250 556929
rect 510284 556895 510318 556929
rect 510352 556895 510386 556929
rect 509493 556784 509527 556818
rect 509493 556716 509527 556750
rect 509493 556648 509527 556682
rect 509493 556580 509527 556614
rect 509493 556512 509527 556546
rect 509493 556444 509527 556478
rect 509493 556376 509527 556410
rect 509493 556308 509527 556342
rect 509493 556240 509527 556274
rect 509493 556172 509527 556206
rect 509493 556104 509527 556138
rect 509493 556036 509527 556070
rect 510463 556784 510497 556818
rect 510463 556716 510497 556750
rect 510463 556648 510497 556682
rect 510463 556580 510497 556614
rect 510463 556512 510497 556546
rect 510463 556444 510497 556478
rect 510463 556376 510497 556410
rect 510463 556308 510497 556342
rect 510463 556240 510497 556274
rect 510463 556172 510497 556206
rect 510463 556104 510497 556138
rect 510463 556036 510497 556070
rect 509604 555925 509638 555959
rect 509672 555925 509706 555959
rect 509740 555925 509774 555959
rect 509808 555925 509842 555959
rect 509876 555925 509910 555959
rect 509944 555925 509978 555959
rect 510012 555925 510046 555959
rect 510080 555925 510114 555959
rect 510148 555925 510182 555959
rect 510216 555925 510250 555959
rect 510284 555925 510318 555959
rect 510352 555925 510386 555959
rect 515450 556895 515484 556929
rect 515518 556895 515552 556929
rect 515586 556895 515620 556929
rect 515654 556895 515688 556929
rect 515722 556895 515756 556929
rect 515790 556895 515824 556929
rect 515858 556895 515892 556929
rect 515926 556895 515960 556929
rect 515994 556895 516028 556929
rect 516062 556895 516096 556929
rect 516130 556895 516164 556929
rect 516198 556895 516232 556929
rect 515339 556784 515373 556818
rect 515339 556716 515373 556750
rect 515339 556648 515373 556682
rect 515339 556580 515373 556614
rect 515339 556512 515373 556546
rect 515339 556444 515373 556478
rect 515339 556376 515373 556410
rect 515339 556308 515373 556342
rect 515339 556240 515373 556274
rect 515339 556172 515373 556206
rect 515339 556104 515373 556138
rect 515339 556036 515373 556070
rect 516309 556784 516343 556818
rect 516309 556716 516343 556750
rect 516309 556648 516343 556682
rect 516309 556580 516343 556614
rect 516309 556512 516343 556546
rect 516309 556444 516343 556478
rect 516309 556376 516343 556410
rect 516309 556308 516343 556342
rect 516309 556240 516343 556274
rect 516309 556172 516343 556206
rect 516309 556104 516343 556138
rect 516309 556036 516343 556070
rect 515450 555925 515484 555959
rect 515518 555925 515552 555959
rect 515586 555925 515620 555959
rect 515654 555925 515688 555959
rect 515722 555925 515756 555959
rect 515790 555925 515824 555959
rect 515858 555925 515892 555959
rect 515926 555925 515960 555959
rect 515994 555925 516028 555959
rect 516062 555925 516096 555959
rect 516130 555925 516164 555959
rect 516198 555925 516232 555959
<< nsubdiffcont >>
rect 509106 557354 509140 557388
rect 509174 557354 509208 557388
rect 509242 557354 509276 557388
rect 509310 557354 509344 557388
rect 509378 557354 509412 557388
rect 509446 557354 509480 557388
rect 509514 557354 509548 557388
rect 509582 557354 509616 557388
rect 509650 557354 509684 557388
rect 509718 557354 509752 557388
rect 509786 557354 509820 557388
rect 509854 557354 509888 557388
rect 509922 557354 509956 557388
rect 509990 557354 510024 557388
rect 510058 557354 510092 557388
rect 510126 557354 510160 557388
rect 510194 557354 510228 557388
rect 510262 557354 510296 557388
rect 510330 557354 510364 557388
rect 510398 557354 510432 557388
rect 510466 557354 510500 557388
rect 510534 557354 510568 557388
rect 510602 557354 510636 557388
rect 510670 557354 510704 557388
rect 510738 557354 510772 557388
rect 510806 557354 510840 557388
rect 510874 557354 510908 557388
rect 509034 557282 509068 557316
rect 509034 557214 509068 557248
rect 509034 557146 509068 557180
rect 509034 557078 509068 557112
rect 509034 557010 509068 557044
rect 509034 556942 509068 556976
rect 510946 557282 510980 557316
rect 510946 557214 510980 557248
rect 510946 557146 510980 557180
rect 510946 557078 510980 557112
rect 510946 557010 510980 557044
rect 510946 556942 510980 556976
rect 509034 556874 509068 556908
rect 509034 556806 509068 556840
rect 509034 556738 509068 556772
rect 509034 556670 509068 556704
rect 509034 556602 509068 556636
rect 509034 556534 509068 556568
rect 509034 556466 509068 556500
rect 509034 556398 509068 556432
rect 509034 556330 509068 556364
rect 509034 556262 509068 556296
rect 509034 556194 509068 556228
rect 509034 556126 509068 556160
rect 509034 556058 509068 556092
rect 509034 555990 509068 556024
rect 509034 555922 509068 555956
rect 510946 556874 510980 556908
rect 510946 556806 510980 556840
rect 510946 556738 510980 556772
rect 510946 556670 510980 556704
rect 510946 556602 510980 556636
rect 510946 556534 510980 556568
rect 510946 556466 510980 556500
rect 510946 556398 510980 556432
rect 510946 556330 510980 556364
rect 510946 556262 510980 556296
rect 510946 556194 510980 556228
rect 510946 556126 510980 556160
rect 510946 556058 510980 556092
rect 510946 555990 510980 556024
rect 509034 555854 509068 555888
rect 509034 555786 509068 555820
rect 509034 555718 509068 555752
rect 509034 555650 509068 555684
rect 509034 555582 509068 555616
rect 509034 555514 509068 555548
rect 510946 555922 510980 555956
rect 510946 555854 510980 555888
rect 510946 555786 510980 555820
rect 510946 555718 510980 555752
rect 510946 555650 510980 555684
rect 510946 555582 510980 555616
rect 510946 555514 510980 555548
rect 509106 555442 509140 555476
rect 509174 555442 509208 555476
rect 509242 555442 509276 555476
rect 509310 555442 509344 555476
rect 509378 555442 509412 555476
rect 509446 555442 509480 555476
rect 509514 555442 509548 555476
rect 509582 555442 509616 555476
rect 509650 555442 509684 555476
rect 509718 555442 509752 555476
rect 509786 555442 509820 555476
rect 509854 555442 509888 555476
rect 509922 555442 509956 555476
rect 509990 555442 510024 555476
rect 510058 555442 510092 555476
rect 510126 555442 510160 555476
rect 510194 555442 510228 555476
rect 510262 555442 510296 555476
rect 510330 555442 510364 555476
rect 510398 555442 510432 555476
rect 510466 555442 510500 555476
rect 510534 555442 510568 555476
rect 510602 555442 510636 555476
rect 510670 555442 510704 555476
rect 510738 555442 510772 555476
rect 510806 555442 510840 555476
rect 510874 555442 510908 555476
rect 514952 557354 514986 557388
rect 515020 557354 515054 557388
rect 515088 557354 515122 557388
rect 515156 557354 515190 557388
rect 515224 557354 515258 557388
rect 515292 557354 515326 557388
rect 515360 557354 515394 557388
rect 515428 557354 515462 557388
rect 515496 557354 515530 557388
rect 515564 557354 515598 557388
rect 515632 557354 515666 557388
rect 515700 557354 515734 557388
rect 515768 557354 515802 557388
rect 515836 557354 515870 557388
rect 515904 557354 515938 557388
rect 515972 557354 516006 557388
rect 516040 557354 516074 557388
rect 516108 557354 516142 557388
rect 516176 557354 516210 557388
rect 516244 557354 516278 557388
rect 516312 557354 516346 557388
rect 516380 557354 516414 557388
rect 516448 557354 516482 557388
rect 516516 557354 516550 557388
rect 516584 557354 516618 557388
rect 516652 557354 516686 557388
rect 516720 557354 516754 557388
rect 514880 557282 514914 557316
rect 514880 557214 514914 557248
rect 514880 557146 514914 557180
rect 514880 557078 514914 557112
rect 514880 557010 514914 557044
rect 514880 556942 514914 556976
rect 516792 557282 516826 557316
rect 516792 557214 516826 557248
rect 516792 557146 516826 557180
rect 516792 557078 516826 557112
rect 516792 557010 516826 557044
rect 516792 556942 516826 556976
rect 514880 556874 514914 556908
rect 514880 556806 514914 556840
rect 514880 556738 514914 556772
rect 514880 556670 514914 556704
rect 514880 556602 514914 556636
rect 514880 556534 514914 556568
rect 514880 556466 514914 556500
rect 514880 556398 514914 556432
rect 514880 556330 514914 556364
rect 514880 556262 514914 556296
rect 514880 556194 514914 556228
rect 514880 556126 514914 556160
rect 514880 556058 514914 556092
rect 514880 555990 514914 556024
rect 514880 555922 514914 555956
rect 516792 556874 516826 556908
rect 516792 556806 516826 556840
rect 516792 556738 516826 556772
rect 516792 556670 516826 556704
rect 516792 556602 516826 556636
rect 516792 556534 516826 556568
rect 516792 556466 516826 556500
rect 516792 556398 516826 556432
rect 516792 556330 516826 556364
rect 516792 556262 516826 556296
rect 516792 556194 516826 556228
rect 516792 556126 516826 556160
rect 516792 556058 516826 556092
rect 516792 555990 516826 556024
rect 514880 555854 514914 555888
rect 514880 555786 514914 555820
rect 514880 555718 514914 555752
rect 514880 555650 514914 555684
rect 514880 555582 514914 555616
rect 514880 555514 514914 555548
rect 516792 555922 516826 555956
rect 516792 555854 516826 555888
rect 516792 555786 516826 555820
rect 516792 555718 516826 555752
rect 516792 555650 516826 555684
rect 516792 555582 516826 555616
rect 516792 555514 516826 555548
rect 514952 555442 514986 555476
rect 515020 555442 515054 555476
rect 515088 555442 515122 555476
rect 515156 555442 515190 555476
rect 515224 555442 515258 555476
rect 515292 555442 515326 555476
rect 515360 555442 515394 555476
rect 515428 555442 515462 555476
rect 515496 555442 515530 555476
rect 515564 555442 515598 555476
rect 515632 555442 515666 555476
rect 515700 555442 515734 555476
rect 515768 555442 515802 555476
rect 515836 555442 515870 555476
rect 515904 555442 515938 555476
rect 515972 555442 516006 555476
rect 516040 555442 516074 555476
rect 516108 555442 516142 555476
rect 516176 555442 516210 555476
rect 516244 555442 516278 555476
rect 516312 555442 516346 555476
rect 516380 555442 516414 555476
rect 516448 555442 516482 555476
rect 516516 555442 516550 555476
rect 516584 555442 516618 555476
rect 516652 555442 516686 555476
rect 516720 555442 516754 555476
<< ndiode >>
rect 509595 558484 510395 558527
rect 509595 557770 509638 558484
rect 510352 557770 510395 558484
rect 509595 557727 510395 557770
rect 515441 558484 516241 558527
rect 515441 557770 515484 558484
rect 516198 557770 516241 558484
rect 515441 557727 516241 557770
rect 509595 556784 510395 556827
rect 509595 556070 509638 556784
rect 510352 556070 510395 556784
rect 509595 556027 510395 556070
rect 515441 556784 516241 556827
rect 515441 556070 515484 556784
rect 516198 556070 516241 556784
rect 515441 556027 516241 556070
<< ndiodec >>
rect 509638 557770 510352 558484
rect 515484 557770 516198 558484
rect 509638 556070 510352 556784
rect 515484 556070 516198 556784
<< locali >>
rect 509567 558703 510417 558715
rect 509567 558629 509615 558703
rect 510369 558629 510417 558703
rect 515413 558703 516263 558715
rect 515413 558629 515461 558703
rect 516215 558629 516263 558703
rect 509493 558595 509604 558629
rect 509638 558595 509672 558597
rect 509706 558595 509740 558597
rect 509774 558595 509808 558597
rect 509842 558595 509876 558597
rect 509910 558595 509944 558597
rect 509978 558595 510012 558597
rect 510046 558595 510080 558597
rect 510114 558595 510148 558597
rect 510182 558595 510216 558597
rect 510250 558595 510284 558597
rect 510318 558595 510352 558597
rect 510386 558595 510497 558629
rect 509493 558518 509527 558595
rect 509567 558585 510417 558595
rect 510463 558518 510497 558595
rect 509493 558450 509527 558484
rect 509493 558382 509527 558416
rect 509493 558314 509527 558348
rect 509493 558246 509527 558280
rect 509493 558178 509527 558212
rect 509493 558110 509527 558144
rect 509493 558042 509527 558076
rect 509493 557974 509527 558008
rect 509493 557906 509527 557940
rect 509493 557838 509527 557872
rect 509493 557770 509527 557804
rect 509591 558504 510399 558515
rect 509591 557750 509618 558504
rect 510372 557750 510399 558504
rect 509591 557739 510399 557750
rect 510463 558450 510497 558484
rect 510463 558382 510497 558416
rect 510463 558314 510497 558348
rect 510463 558246 510497 558280
rect 510463 558178 510497 558212
rect 510463 558110 510497 558144
rect 510463 558042 510497 558076
rect 510463 557974 510497 558008
rect 510463 557906 510497 557940
rect 510463 557838 510497 557872
rect 510463 557770 510497 557804
rect 509493 557659 509527 557736
rect 510463 557659 510497 557736
rect 509493 557625 509604 557659
rect 509638 557625 509672 557659
rect 509706 557625 509740 557659
rect 509774 557625 509808 557659
rect 509842 557625 509876 557659
rect 509910 557625 509944 557659
rect 509978 557625 510012 557659
rect 510046 557625 510080 557659
rect 510114 557625 510148 557659
rect 510182 557625 510216 557659
rect 510250 557625 510284 557659
rect 510318 557625 510352 557659
rect 510386 557625 510497 557659
rect 515339 558595 515450 558629
rect 515484 558595 515518 558597
rect 515552 558595 515586 558597
rect 515620 558595 515654 558597
rect 515688 558595 515722 558597
rect 515756 558595 515790 558597
rect 515824 558595 515858 558597
rect 515892 558595 515926 558597
rect 515960 558595 515994 558597
rect 516028 558595 516062 558597
rect 516096 558595 516130 558597
rect 516164 558595 516198 558597
rect 516232 558595 516343 558629
rect 515339 558518 515373 558595
rect 515413 558585 516263 558595
rect 516309 558518 516343 558595
rect 515339 558450 515373 558484
rect 515339 558382 515373 558416
rect 515339 558314 515373 558348
rect 515339 558246 515373 558280
rect 515339 558178 515373 558212
rect 515339 558110 515373 558144
rect 515339 558042 515373 558076
rect 515339 557974 515373 558008
rect 515339 557906 515373 557940
rect 515339 557838 515373 557872
rect 515339 557770 515373 557804
rect 515437 558504 516245 558515
rect 515437 557750 515464 558504
rect 516218 557750 516245 558504
rect 515437 557739 516245 557750
rect 516309 558450 516343 558484
rect 516309 558382 516343 558416
rect 516309 558314 516343 558348
rect 516309 558246 516343 558280
rect 516309 558178 516343 558212
rect 516309 558110 516343 558144
rect 516309 558042 516343 558076
rect 516309 557974 516343 558008
rect 516309 557906 516343 557940
rect 516309 557838 516343 557872
rect 516309 557770 516343 557804
rect 515339 557659 515373 557736
rect 516309 557659 516343 557736
rect 515339 557625 515450 557659
rect 515484 557625 515518 557659
rect 515552 557625 515586 557659
rect 515620 557625 515654 557659
rect 515688 557625 515722 557659
rect 515756 557625 515790 557659
rect 515824 557625 515858 557659
rect 515892 557625 515926 557659
rect 515960 557625 515994 557659
rect 516028 557625 516062 557659
rect 516096 557625 516130 557659
rect 516164 557625 516198 557659
rect 516232 557625 516343 557659
rect 509034 557354 509106 557388
rect 509140 557354 509174 557388
rect 509208 557354 509242 557388
rect 509276 557354 509310 557388
rect 509344 557354 509378 557388
rect 509412 557354 509446 557388
rect 509480 557354 509514 557388
rect 509548 557354 509582 557388
rect 509616 557354 509650 557388
rect 509684 557354 509718 557388
rect 509752 557354 509786 557388
rect 509820 557354 509854 557388
rect 509888 557354 509922 557388
rect 509956 557354 509990 557388
rect 510024 557354 510058 557388
rect 510092 557354 510126 557388
rect 510160 557354 510194 557388
rect 510228 557354 510262 557388
rect 510296 557354 510330 557388
rect 510364 557354 510398 557388
rect 510432 557354 510466 557388
rect 510500 557354 510534 557388
rect 510568 557354 510602 557388
rect 510636 557354 510670 557388
rect 510704 557354 510738 557388
rect 510772 557354 510806 557388
rect 510840 557354 510874 557388
rect 510908 557354 510980 557388
rect 509034 557316 509068 557354
rect 509034 557248 509068 557282
rect 509034 557180 509068 557214
rect 509034 557112 509068 557146
rect 509034 557044 509068 557078
rect 509034 556976 509068 557010
rect 510946 557316 510980 557354
rect 510946 557248 510980 557282
rect 510946 557180 510980 557214
rect 510946 557112 510980 557146
rect 510946 557044 510980 557078
rect 509034 556908 509068 556942
rect 509577 556952 510407 556985
rect 509577 556929 509615 556952
rect 509649 556929 509687 556952
rect 509721 556929 509759 556952
rect 509793 556929 509831 556952
rect 509865 556929 509903 556952
rect 509937 556929 509975 556952
rect 510009 556929 510047 556952
rect 510081 556929 510119 556952
rect 510153 556929 510191 556952
rect 510225 556929 510263 556952
rect 510297 556929 510335 556952
rect 510369 556929 510407 556952
rect 510946 556976 510980 557010
rect 509034 556840 509068 556874
rect 509034 556772 509068 556806
rect 509034 556704 509068 556738
rect 509034 556636 509068 556670
rect 509034 556568 509068 556602
rect 509034 556500 509068 556534
rect 509034 556432 509068 556466
rect 509034 556364 509068 556398
rect 509034 556296 509068 556330
rect 509034 556228 509068 556262
rect 509034 556160 509068 556194
rect 509034 556092 509068 556126
rect 509034 556024 509068 556058
rect 509034 555956 509068 555990
rect 509493 556895 509604 556929
rect 509649 556918 509672 556929
rect 509721 556918 509740 556929
rect 509793 556918 509808 556929
rect 509865 556918 509876 556929
rect 509937 556918 509944 556929
rect 510009 556918 510012 556929
rect 509638 556895 509672 556918
rect 509706 556895 509740 556918
rect 509774 556895 509808 556918
rect 509842 556895 509876 556918
rect 509910 556895 509944 556918
rect 509978 556895 510012 556918
rect 510046 556918 510047 556929
rect 510114 556918 510119 556929
rect 510182 556918 510191 556929
rect 510250 556918 510263 556929
rect 510318 556918 510335 556929
rect 510046 556895 510080 556918
rect 510114 556895 510148 556918
rect 510182 556895 510216 556918
rect 510250 556895 510284 556918
rect 510318 556895 510352 556918
rect 510386 556895 510497 556929
rect 509493 556818 509527 556895
rect 509577 556885 510407 556895
rect 510463 556818 510497 556895
rect 509493 556750 509527 556784
rect 509493 556682 509527 556716
rect 509493 556614 509527 556648
rect 509493 556546 509527 556580
rect 509493 556478 509527 556512
rect 509493 556410 509527 556444
rect 509493 556342 509527 556376
rect 509493 556274 509527 556308
rect 509493 556206 509527 556240
rect 509493 556138 509527 556172
rect 509493 556070 509527 556104
rect 509591 556804 510399 556815
rect 509591 556050 509618 556804
rect 510372 556050 510399 556804
rect 509591 556039 510399 556050
rect 510463 556750 510497 556784
rect 510463 556682 510497 556716
rect 510463 556614 510497 556648
rect 510463 556546 510497 556580
rect 510463 556478 510497 556512
rect 510463 556410 510497 556444
rect 510463 556342 510497 556376
rect 510463 556274 510497 556308
rect 510463 556206 510497 556240
rect 510463 556138 510497 556172
rect 510463 556070 510497 556104
rect 509493 555959 509527 556036
rect 510463 555959 510497 556036
rect 509493 555925 509604 555959
rect 509638 555925 509672 555959
rect 509706 555925 509740 555959
rect 509774 555925 509808 555959
rect 509842 555925 509876 555959
rect 509910 555925 509944 555959
rect 509978 555925 510012 555959
rect 510046 555925 510080 555959
rect 510114 555925 510148 555959
rect 510182 555925 510216 555959
rect 510250 555925 510284 555959
rect 510318 555925 510352 555959
rect 510386 555925 510497 555959
rect 510946 556908 510980 556942
rect 510946 556840 510980 556874
rect 510946 556772 510980 556806
rect 510946 556704 510980 556738
rect 510946 556636 510980 556670
rect 510946 556568 510980 556602
rect 510946 556500 510980 556534
rect 510946 556432 510980 556466
rect 510946 556364 510980 556398
rect 510946 556296 510980 556330
rect 510946 556228 510980 556262
rect 510946 556160 510980 556194
rect 510946 556092 510980 556126
rect 510946 556024 510980 556058
rect 510946 555956 510980 555990
rect 509034 555888 509068 555922
rect 509034 555820 509068 555854
rect 509034 555752 509068 555786
rect 509034 555684 509068 555718
rect 509034 555616 509068 555650
rect 509034 555548 509068 555582
rect 509034 555476 509068 555514
rect 510946 555888 510980 555922
rect 510946 555820 510980 555854
rect 510946 555752 510980 555786
rect 510946 555684 510980 555718
rect 510946 555616 510980 555650
rect 510946 555548 510980 555582
rect 510946 555476 510980 555514
rect 509034 555442 509106 555476
rect 509140 555442 509174 555476
rect 509208 555442 509242 555476
rect 509276 555442 509310 555476
rect 509344 555442 509378 555476
rect 509412 555442 509446 555476
rect 509480 555442 509514 555476
rect 509548 555442 509582 555476
rect 509616 555442 509650 555476
rect 509684 555442 509718 555476
rect 509752 555442 509786 555476
rect 509820 555442 509854 555476
rect 509888 555442 509922 555476
rect 509956 555442 509990 555476
rect 510024 555442 510058 555476
rect 510092 555442 510126 555476
rect 510160 555442 510194 555476
rect 510228 555442 510262 555476
rect 510296 555442 510330 555476
rect 510364 555442 510398 555476
rect 510432 555442 510466 555476
rect 510500 555442 510534 555476
rect 510568 555442 510602 555476
rect 510636 555442 510670 555476
rect 510704 555442 510738 555476
rect 510772 555442 510806 555476
rect 510840 555442 510874 555476
rect 510908 555442 510980 555476
rect 514880 557354 514952 557388
rect 514986 557354 515020 557388
rect 515054 557354 515088 557388
rect 515122 557354 515156 557388
rect 515190 557354 515224 557388
rect 515258 557354 515292 557388
rect 515326 557354 515360 557388
rect 515394 557354 515428 557388
rect 515462 557354 515496 557388
rect 515530 557354 515564 557388
rect 515598 557354 515632 557388
rect 515666 557354 515700 557388
rect 515734 557354 515768 557388
rect 515802 557354 515836 557388
rect 515870 557354 515904 557388
rect 515938 557354 515972 557388
rect 516006 557354 516040 557388
rect 516074 557354 516108 557388
rect 516142 557354 516176 557388
rect 516210 557354 516244 557388
rect 516278 557354 516312 557388
rect 516346 557354 516380 557388
rect 516414 557354 516448 557388
rect 516482 557354 516516 557388
rect 516550 557354 516584 557388
rect 516618 557354 516652 557388
rect 516686 557354 516720 557388
rect 516754 557354 516826 557388
rect 514880 557316 514914 557354
rect 514880 557248 514914 557282
rect 514880 557180 514914 557214
rect 514880 557112 514914 557146
rect 514880 557044 514914 557078
rect 514880 556976 514914 557010
rect 516792 557316 516826 557354
rect 516792 557248 516826 557282
rect 516792 557180 516826 557214
rect 516792 557112 516826 557146
rect 516792 557044 516826 557078
rect 514880 556908 514914 556942
rect 515423 556952 516253 556985
rect 515423 556929 515461 556952
rect 515495 556929 515533 556952
rect 515567 556929 515605 556952
rect 515639 556929 515677 556952
rect 515711 556929 515749 556952
rect 515783 556929 515821 556952
rect 515855 556929 515893 556952
rect 515927 556929 515965 556952
rect 515999 556929 516037 556952
rect 516071 556929 516109 556952
rect 516143 556929 516181 556952
rect 516215 556929 516253 556952
rect 516792 556976 516826 557010
rect 514880 556840 514914 556874
rect 514880 556772 514914 556806
rect 514880 556704 514914 556738
rect 514880 556636 514914 556670
rect 514880 556568 514914 556602
rect 514880 556500 514914 556534
rect 514880 556432 514914 556466
rect 514880 556364 514914 556398
rect 514880 556296 514914 556330
rect 514880 556228 514914 556262
rect 514880 556160 514914 556194
rect 514880 556092 514914 556126
rect 514880 556024 514914 556058
rect 514880 555956 514914 555990
rect 515339 556895 515450 556929
rect 515495 556918 515518 556929
rect 515567 556918 515586 556929
rect 515639 556918 515654 556929
rect 515711 556918 515722 556929
rect 515783 556918 515790 556929
rect 515855 556918 515858 556929
rect 515484 556895 515518 556918
rect 515552 556895 515586 556918
rect 515620 556895 515654 556918
rect 515688 556895 515722 556918
rect 515756 556895 515790 556918
rect 515824 556895 515858 556918
rect 515892 556918 515893 556929
rect 515960 556918 515965 556929
rect 516028 556918 516037 556929
rect 516096 556918 516109 556929
rect 516164 556918 516181 556929
rect 515892 556895 515926 556918
rect 515960 556895 515994 556918
rect 516028 556895 516062 556918
rect 516096 556895 516130 556918
rect 516164 556895 516198 556918
rect 516232 556895 516343 556929
rect 515339 556818 515373 556895
rect 515423 556885 516253 556895
rect 516309 556818 516343 556895
rect 515339 556750 515373 556784
rect 515339 556682 515373 556716
rect 515339 556614 515373 556648
rect 515339 556546 515373 556580
rect 515339 556478 515373 556512
rect 515339 556410 515373 556444
rect 515339 556342 515373 556376
rect 515339 556274 515373 556308
rect 515339 556206 515373 556240
rect 515339 556138 515373 556172
rect 515339 556070 515373 556104
rect 515437 556804 516245 556815
rect 515437 556050 515464 556804
rect 516218 556050 516245 556804
rect 515437 556039 516245 556050
rect 516309 556750 516343 556784
rect 516309 556682 516343 556716
rect 516309 556614 516343 556648
rect 516309 556546 516343 556580
rect 516309 556478 516343 556512
rect 516309 556410 516343 556444
rect 516309 556342 516343 556376
rect 516309 556274 516343 556308
rect 516309 556206 516343 556240
rect 516309 556138 516343 556172
rect 516309 556070 516343 556104
rect 515339 555959 515373 556036
rect 516309 555959 516343 556036
rect 515339 555925 515450 555959
rect 515484 555925 515518 555959
rect 515552 555925 515586 555959
rect 515620 555925 515654 555959
rect 515688 555925 515722 555959
rect 515756 555925 515790 555959
rect 515824 555925 515858 555959
rect 515892 555925 515926 555959
rect 515960 555925 515994 555959
rect 516028 555925 516062 555959
rect 516096 555925 516130 555959
rect 516164 555925 516198 555959
rect 516232 555925 516343 555959
rect 516792 556908 516826 556942
rect 516792 556840 516826 556874
rect 516792 556772 516826 556806
rect 516792 556704 516826 556738
rect 516792 556636 516826 556670
rect 516792 556568 516826 556602
rect 516792 556500 516826 556534
rect 516792 556432 516826 556466
rect 516792 556364 516826 556398
rect 516792 556296 516826 556330
rect 516792 556228 516826 556262
rect 516792 556160 516826 556194
rect 516792 556092 516826 556126
rect 516792 556024 516826 556058
rect 516792 555956 516826 555990
rect 514880 555888 514914 555922
rect 514880 555820 514914 555854
rect 514880 555752 514914 555786
rect 514880 555684 514914 555718
rect 514880 555616 514914 555650
rect 514880 555548 514914 555582
rect 514880 555476 514914 555514
rect 516792 555888 516826 555922
rect 516792 555820 516826 555854
rect 516792 555752 516826 555786
rect 516792 555684 516826 555718
rect 516792 555616 516826 555650
rect 516792 555548 516826 555582
rect 516792 555476 516826 555514
rect 514880 555442 514952 555476
rect 514986 555442 515020 555476
rect 515054 555442 515088 555476
rect 515122 555442 515156 555476
rect 515190 555442 515224 555476
rect 515258 555442 515292 555476
rect 515326 555442 515360 555476
rect 515394 555442 515428 555476
rect 515462 555442 515496 555476
rect 515530 555442 515564 555476
rect 515598 555442 515632 555476
rect 515666 555442 515700 555476
rect 515734 555442 515768 555476
rect 515802 555442 515836 555476
rect 515870 555442 515904 555476
rect 515938 555442 515972 555476
rect 516006 555442 516040 555476
rect 516074 555442 516108 555476
rect 516142 555442 516176 555476
rect 516210 555442 516244 555476
rect 516278 555442 516312 555476
rect 516346 555442 516380 555476
rect 516414 555442 516448 555476
rect 516482 555442 516516 555476
rect 516550 555442 516584 555476
rect 516618 555442 516652 555476
rect 516686 555442 516720 555476
rect 516754 555442 516826 555476
<< viali >>
rect 509615 558629 510369 558703
rect 515461 558629 516215 558703
rect 509615 558597 509638 558629
rect 509638 558597 509672 558629
rect 509672 558597 509706 558629
rect 509706 558597 509740 558629
rect 509740 558597 509774 558629
rect 509774 558597 509808 558629
rect 509808 558597 509842 558629
rect 509842 558597 509876 558629
rect 509876 558597 509910 558629
rect 509910 558597 509944 558629
rect 509944 558597 509978 558629
rect 509978 558597 510012 558629
rect 510012 558597 510046 558629
rect 510046 558597 510080 558629
rect 510080 558597 510114 558629
rect 510114 558597 510148 558629
rect 510148 558597 510182 558629
rect 510182 558597 510216 558629
rect 510216 558597 510250 558629
rect 510250 558597 510284 558629
rect 510284 558597 510318 558629
rect 510318 558597 510352 558629
rect 510352 558597 510369 558629
rect 509618 558484 510372 558504
rect 509618 557770 509638 558484
rect 509638 557770 510352 558484
rect 510352 557770 510372 558484
rect 509618 557750 510372 557770
rect 515461 558597 515484 558629
rect 515484 558597 515518 558629
rect 515518 558597 515552 558629
rect 515552 558597 515586 558629
rect 515586 558597 515620 558629
rect 515620 558597 515654 558629
rect 515654 558597 515688 558629
rect 515688 558597 515722 558629
rect 515722 558597 515756 558629
rect 515756 558597 515790 558629
rect 515790 558597 515824 558629
rect 515824 558597 515858 558629
rect 515858 558597 515892 558629
rect 515892 558597 515926 558629
rect 515926 558597 515960 558629
rect 515960 558597 515994 558629
rect 515994 558597 516028 558629
rect 516028 558597 516062 558629
rect 516062 558597 516096 558629
rect 516096 558597 516130 558629
rect 516130 558597 516164 558629
rect 516164 558597 516198 558629
rect 516198 558597 516215 558629
rect 515464 558484 516218 558504
rect 515464 557770 515484 558484
rect 515484 557770 516198 558484
rect 516198 557770 516218 558484
rect 515464 557750 516218 557770
rect 509615 556929 509649 556952
rect 509687 556929 509721 556952
rect 509759 556929 509793 556952
rect 509831 556929 509865 556952
rect 509903 556929 509937 556952
rect 509975 556929 510009 556952
rect 510047 556929 510081 556952
rect 510119 556929 510153 556952
rect 510191 556929 510225 556952
rect 510263 556929 510297 556952
rect 510335 556929 510369 556952
rect 509615 556918 509638 556929
rect 509638 556918 509649 556929
rect 509687 556918 509706 556929
rect 509706 556918 509721 556929
rect 509759 556918 509774 556929
rect 509774 556918 509793 556929
rect 509831 556918 509842 556929
rect 509842 556918 509865 556929
rect 509903 556918 509910 556929
rect 509910 556918 509937 556929
rect 509975 556918 509978 556929
rect 509978 556918 510009 556929
rect 510047 556918 510080 556929
rect 510080 556918 510081 556929
rect 510119 556918 510148 556929
rect 510148 556918 510153 556929
rect 510191 556918 510216 556929
rect 510216 556918 510225 556929
rect 510263 556918 510284 556929
rect 510284 556918 510297 556929
rect 510335 556918 510352 556929
rect 510352 556918 510369 556929
rect 509618 556784 510372 556804
rect 509618 556070 509638 556784
rect 509638 556070 510352 556784
rect 510352 556070 510372 556784
rect 509618 556050 510372 556070
rect 515461 556929 515495 556952
rect 515533 556929 515567 556952
rect 515605 556929 515639 556952
rect 515677 556929 515711 556952
rect 515749 556929 515783 556952
rect 515821 556929 515855 556952
rect 515893 556929 515927 556952
rect 515965 556929 515999 556952
rect 516037 556929 516071 556952
rect 516109 556929 516143 556952
rect 516181 556929 516215 556952
rect 515461 556918 515484 556929
rect 515484 556918 515495 556929
rect 515533 556918 515552 556929
rect 515552 556918 515567 556929
rect 515605 556918 515620 556929
rect 515620 556918 515639 556929
rect 515677 556918 515688 556929
rect 515688 556918 515711 556929
rect 515749 556918 515756 556929
rect 515756 556918 515783 556929
rect 515821 556918 515824 556929
rect 515824 556918 515855 556929
rect 515893 556918 515926 556929
rect 515926 556918 515927 556929
rect 515965 556918 515994 556929
rect 515994 556918 515999 556929
rect 516037 556918 516062 556929
rect 516062 556918 516071 556929
rect 516109 556918 516130 556929
rect 516130 556918 516143 556929
rect 516181 556918 516198 556929
rect 516198 556918 516215 556929
rect 515464 556784 516218 556804
rect 515464 556070 515484 556784
rect 515484 556070 516198 556784
rect 516198 556070 516218 556784
rect 515464 556050 516218 556070
<< metal1 >>
rect 7832 687526 9320 688392
rect 11747 687437 13958 688451
rect 7832 684278 9320 685144
rect 11747 684228 13958 685242
rect 509563 558703 510429 560138
rect 509563 558650 509615 558703
rect 509567 558597 509615 558650
rect 510369 558650 510429 558703
rect 515408 558703 516274 560138
rect 515408 558650 515461 558703
rect 510369 558597 510417 558650
rect 509567 558585 510417 558597
rect 515413 558597 515461 558650
rect 516215 558650 516274 558703
rect 516215 558597 516263 558650
rect 515413 558585 516263 558597
rect 509577 558504 510407 558525
rect 509577 557750 509618 558504
rect 510372 557750 510407 558504
rect 509577 556952 510407 557750
rect 509577 556918 509615 556952
rect 509649 556918 509687 556952
rect 509721 556918 509759 556952
rect 509793 556918 509831 556952
rect 509865 556918 509903 556952
rect 509937 556918 509975 556952
rect 510009 556918 510047 556952
rect 510081 556918 510119 556952
rect 510153 556918 510191 556952
rect 510225 556918 510263 556952
rect 510297 556918 510335 556952
rect 510369 556918 510407 556952
rect 509577 556885 510407 556918
rect 515423 558504 516253 558525
rect 515423 557750 515464 558504
rect 516218 557750 516253 558504
rect 515423 556952 516253 557750
rect 515423 556918 515461 556952
rect 515495 556918 515533 556952
rect 515567 556918 515605 556952
rect 515639 556918 515677 556952
rect 515711 556918 515749 556952
rect 515783 556918 515821 556952
rect 515855 556918 515893 556952
rect 515927 556918 515965 556952
rect 515999 556918 516037 556952
rect 516071 556918 516109 556952
rect 516143 556918 516181 556952
rect 516215 556918 516253 556952
rect 515423 556885 516253 556918
rect 509587 556804 510407 556825
rect 509587 556223 509618 556804
rect 509465 556050 509618 556223
rect 510372 556223 510407 556804
rect 515433 556804 516253 556825
rect 515433 556223 515464 556804
rect 510372 556050 510479 556223
rect 509465 554012 510479 556050
rect 515349 556050 515464 556223
rect 516218 556223 516253 556804
rect 516218 556050 516363 556223
rect 515349 554012 516363 556050
rect 526048 510660 526648 597175
rect 63230 491883 63600 494452
rect 65030 491868 65400 494488
rect 526262 442316 526402 500309
rect 471628 442176 526402 442316
rect 482380 415325 482520 417119
rect 482380 415185 506016 415325
<< metal2 >>
rect 7839 556625 8839 689046
rect 9331 687494 10976 688497
rect 9712 682286 10565 685179
rect 12921 640645 13921 689119
rect 513761 561484 513901 626662
rect 526048 596807 526648 649835
rect 511518 560556 513901 561484
rect 511518 558258 512166 560556
rect 509304 557405 512166 558258
rect 513426 557889 513905 558713
rect 515229 557889 516232 558639
rect 513426 556994 516232 557889
rect 63205 493421 63621 494440
rect 65007 493421 65423 494440
rect 513761 453101 513901 556994
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 17970 688488 18970 702300
rect 9326 687488 18970 688488
rect 510594 688389 525394 702340
rect 566594 702300 571594 704800
rect 568823 693469 569423 702300
rect 17970 685964 18970 687488
rect -800 683292 1700 685242
rect 17970 684964 49842 685964
rect -800 682292 47346 683292
rect -800 680242 1700 682292
rect -800 643842 8110 648642
rect 1660 641850 8110 643842
rect 1660 640850 44988 641850
rect 1660 638642 8110 640850
rect -800 633842 8110 638642
rect 1660 633838 8110 633842
rect -800 564241 1660 564242
rect -800 559442 6373 564241
rect 1573 557634 6373 559442
rect 1573 556634 42612 557634
rect 1573 554242 6373 556634
rect -800 549442 6373 554242
rect 1573 549401 6373 549442
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 39148 506914
rect -800 505620 480 505732
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 38368 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 37420 420470
rect -800 419176 480 419288
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 36524 377248
rect -800 375954 480 376066
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 35440 334026
rect -800 332732 480 332844
rect 35328 324960 35440 333914
rect 36412 325894 36524 377136
rect 37308 326894 37420 420358
rect 38256 327788 38368 464762
rect 39036 328608 39148 506802
rect 41612 481627 42612 556634
rect 43988 484504 44988 640850
rect 46346 494424 47346 682292
rect 48842 496562 49842 684964
rect 568822 684288 569422 693469
rect 526049 683688 569422 684288
rect 526049 664561 526649 683688
rect 582300 680654 584800 682984
rect 568807 680514 584800 680654
rect 526048 649115 526648 664561
rect 568807 626662 568947 680514
rect 582300 677984 584800 680514
rect 582340 639784 584800 644584
rect 582340 629784 584800 634584
rect 513761 626522 568947 626662
rect 583520 589472 584800 589584
rect 517596 588402 583520 588406
rect 517596 588290 584800 588402
rect 517596 588286 583520 588290
rect 48842 495562 65650 496562
rect 46346 493424 63665 494424
rect 64650 493400 65650 495562
rect 41612 480627 45885 481627
rect 513761 415325 513901 453101
rect 505784 415185 513901 415325
rect 452088 374795 452288 374817
tri 452088 332526 452090 374795 ne
rect 452090 363324 452288 374795
rect 454892 374692 455012 374795
tri 454892 366099 454893 374692 ne
rect 454893 366183 455012 374692
tri 455012 366183 455013 374692 sw
tri 452288 363324 452289 366099 sw
rect 53513 328608 53625 331267
rect 39036 328496 53625 328608
rect 55282 327788 55394 331351
rect 38256 327676 55394 327788
rect 57045 326894 57157 331312
rect 37308 326782 57157 326894
rect 58816 325894 58928 331287
rect 36412 325782 58928 325894
rect 60584 324960 60696 331292
rect 35328 324848 60696 324960
rect 62355 323944 62467 331259
rect 16038 323832 62467 323944
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect 16038 290804 16150 323832
rect 64125 322768 64237 331307
rect -800 290692 16150 290804
rect 17454 322656 64237 322768
rect -800 289510 480 289622
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect 17454 247782 17566 322656
rect 65887 321532 65999 331276
rect -800 247670 17566 247782
rect 18914 321420 65999 321532
rect -800 246488 480 246600
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect 18914 120160 19026 321420
rect 67654 320172 67766 331275
rect -800 120048 19026 120160
rect 20370 320060 67766 320172
rect -800 118866 480 118978
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect 20370 76938 20482 320060
rect 69426 318598 69538 331291
rect -800 76826 20482 76938
rect 21956 318486 69538 318598
rect -800 75644 480 75756
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect 21956 33716 22068 318486
rect 71192 317174 71304 331275
rect 452090 331259 452289 363324
rect 454893 365891 455013 366183
rect 457653 366011 457773 374805
rect 460412 369241 460532 374784
rect 463173 372251 463293 374781
rect 465934 374304 466054 374812
rect 517596 374304 517716 588286
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 568389 550562 584800 555362
rect 568389 545362 582340 550562
rect 568389 540562 584800 545362
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 465934 374184 517716 374304
rect 521208 497798 583520 497802
rect 521208 497686 584800 497798
rect 521208 497682 583520 497686
rect 521208 372251 521328 497682
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 463173 372131 521328 372251
rect 524948 453376 583520 453380
rect 524948 453264 584800 453376
rect 524948 453260 583520 453264
rect 524948 369241 525068 453260
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 460412 369121 525068 369241
rect 528935 408954 583520 408957
rect 528935 408842 584800 408954
rect 528935 408837 583520 408842
rect 528935 366011 529055 408837
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 457653 365891 529055 366011
tri 454893 362417 454894 365891 ne
rect 454894 362537 455013 365891
tri 455013 362537 455014 365891 sw
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 454894 362532 583520 362537
rect 454894 362420 584800 362532
rect 454894 362417 583520 362420
rect -800 33604 22068 33716
rect 23136 317062 71304 317174
rect -800 32422 480 32534
rect -800 16910 480 17022
rect -800 15728 480 15840
rect -800 14546 480 14658
rect -800 13364 480 13476
rect 23136 12294 23248 317062
rect 72963 315516 73075 331258
rect -800 12182 23248 12294
rect 24772 315404 73075 315516
rect -800 11000 480 11112
rect -800 9818 480 9930
rect 24772 8748 24884 315404
rect 74729 314070 74841 331259
tri 452090 320998 452091 331259 ne
rect 452091 317354 452289 331259
tri 452289 317354 452291 362417 sw
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 452091 317310 583523 317354
rect 452091 317198 584800 317310
rect 452091 317154 583523 317198
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect -800 8636 24884 8748
rect 26916 313958 74841 314070
rect -800 7454 480 7566
rect -800 6272 480 6384
rect -800 5090 480 5202
rect 26916 4020 27028 313958
rect 583520 313652 584800 313764
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 583520 16910 584800 17022
rect 583520 15728 584800 15840
rect 583520 14546 584800 14658
rect 583520 13364 584800 13476
rect 583520 12182 584800 12294
rect 583520 11000 584800 11112
rect 583520 9818 584800 9930
rect 583520 8636 584800 8748
rect 583520 7454 584800 7566
rect 583520 6272 584800 6384
rect 583520 5090 584800 5202
rect -800 3908 27028 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 510594 688389 525394 702340
rect 495764 552400 582340 555889
rect 495764 550400 496723 552400
rect 498723 550400 499723 552400
rect 501723 550400 502723 552400
rect 504723 550400 505723 552400
rect 507723 550400 508723 552400
rect 510723 550400 511723 552400
rect 513723 550400 514723 552400
rect 516723 550400 517723 552400
rect 519723 550400 582340 552400
rect 495764 549400 582340 550400
rect 495764 547400 496723 549400
rect 498723 547400 499723 549400
rect 501723 547400 502723 549400
rect 504723 547400 505723 549400
rect 507723 547400 508723 549400
rect 510723 547400 511723 549400
rect 513723 547400 514723 549400
rect 516723 547400 517723 549400
rect 519723 547400 582340 549400
rect 495764 546400 582340 547400
rect 495764 544400 496723 546400
rect 498723 544400 499723 546400
rect 501723 544400 502723 546400
rect 504723 544400 505723 546400
rect 507723 544400 508723 546400
rect 510723 544400 511723 546400
rect 513723 544400 514723 546400
rect 516723 544400 517723 546400
rect 519723 544400 582340 546400
rect 495764 543400 582340 544400
rect 495764 541400 496723 543400
rect 498723 541400 499723 543400
rect 501723 541400 502723 543400
rect 504723 541400 505723 543400
rect 507723 541400 508723 543400
rect 510723 541400 511723 543400
rect 513723 541400 514723 543400
rect 516723 541400 517723 543400
rect 519723 541400 582340 543400
rect 495764 541089 582340 541400
rect 495764 540400 528966 541089
rect 495764 538400 496723 540400
rect 498723 538400 499723 540400
rect 501723 538400 502723 540400
rect 504723 538400 505723 540400
rect 507723 538400 508723 540400
rect 510723 538400 511723 540400
rect 513723 538400 514723 540400
rect 516723 538400 517723 540400
rect 519723 538400 528966 540400
rect 495764 537400 528966 538400
rect 495764 535400 496723 537400
rect 498723 535400 499723 537400
rect 501723 535400 502723 537400
rect 504723 535400 505723 537400
rect 507723 535400 508723 537400
rect 510723 535400 511723 537400
rect 513723 535400 514723 537400
rect 516723 535400 517723 537400
rect 519723 535400 528966 537400
rect 495764 534400 528966 535400
rect 495764 532400 496723 534400
rect 498723 532400 499723 534400
rect 501723 532400 502723 534400
rect 504723 532400 505723 534400
rect 507723 532400 508723 534400
rect 510723 532400 511723 534400
rect 513723 532400 514723 534400
rect 516723 532400 517723 534400
rect 519723 532400 528966 534400
rect 495764 531400 528966 532400
rect 495764 529400 496723 531400
rect 498723 529400 499723 531400
rect 501723 529400 502723 531400
rect 504723 529400 505723 531400
rect 507723 529400 508723 531400
rect 510723 529400 511723 531400
rect 513723 529400 514723 531400
rect 516723 529400 517723 531400
rect 519723 529400 528966 531400
rect 495764 528400 528966 529400
rect 495764 526400 496723 528400
rect 498723 526400 499723 528400
rect 501723 526400 502723 528400
rect 504723 526400 505723 528400
rect 507723 526400 508723 528400
rect 510723 526400 511723 528400
rect 513723 526400 514723 528400
rect 516723 526400 517723 528400
rect 519723 526400 528966 528400
rect 495764 525400 528966 526400
rect 495764 523400 496723 525400
rect 498723 523400 499723 525400
rect 501723 523400 502723 525400
rect 504723 523400 505723 525400
rect 507723 523400 508723 525400
rect 510723 523400 511723 525400
rect 513723 523400 514723 525400
rect 516723 523400 517723 525400
rect 519723 523400 528966 525400
rect 495764 522400 528966 523400
rect 495764 520400 496723 522400
rect 498723 520400 499723 522400
rect 501723 520400 502723 522400
rect 504723 520400 505723 522400
rect 507723 520400 508723 522400
rect 510723 520400 511723 522400
rect 513723 520400 514723 522400
rect 516723 520400 517723 522400
rect 519723 520400 528966 522400
rect 495764 519400 528966 520400
rect 495764 517400 496723 519400
rect 498723 517400 499723 519400
rect 501723 517400 502723 519400
rect 504723 517400 505723 519400
rect 507723 517400 508723 519400
rect 510723 517400 511723 519400
rect 513723 517400 514723 519400
rect 516723 517400 517723 519400
rect 519723 517400 528966 519400
rect 495764 516400 528966 517400
rect 495764 514400 496723 516400
rect 498723 514400 499723 516400
rect 501723 514400 502723 516400
rect 504723 514400 505723 516400
rect 507723 514400 508723 516400
rect 510723 514400 511723 516400
rect 513723 514400 514723 516400
rect 516723 514400 517723 516400
rect 519723 514400 528966 516400
rect 495764 513400 528966 514400
rect 495764 511400 496723 513400
rect 498723 511400 499723 513400
rect 501723 511400 502723 513400
rect 504723 511400 505723 513400
rect 507723 511400 508723 513400
rect 510723 511400 511723 513400
rect 513723 511400 514723 513400
rect 516723 511400 517723 513400
rect 519723 511400 528966 513400
rect 495764 511240 528966 511400
rect 495764 510400 524273 511240
rect 528170 510979 528966 511240
rect 495764 508400 496723 510400
rect 498723 508400 499723 510400
rect 501723 508400 502723 510400
rect 504723 508400 505723 510400
rect 507723 508400 508723 510400
rect 510723 508400 511723 510400
rect 513723 508400 514723 510400
rect 516723 508400 517723 510400
rect 519723 508400 524273 510400
rect 528236 510282 528966 510979
rect 495764 507400 524273 508400
rect 495764 505400 496723 507400
rect 498723 505400 499723 507400
rect 501723 505400 502723 507400
rect 504723 505400 505723 507400
rect 507723 505400 508723 507400
rect 510723 505400 511723 507400
rect 513723 505400 514723 507400
rect 516723 505400 517723 507400
rect 519723 505400 524273 507400
rect 495764 504400 524273 505400
rect 495764 502400 496723 504400
rect 498723 502400 499723 504400
rect 501723 502400 502723 504400
rect 504723 502400 505723 504400
rect 507723 502400 508723 504400
rect 510723 502400 511723 504400
rect 513723 502400 514723 504400
rect 516723 502400 517723 504400
rect 519723 502400 524273 504400
rect 495764 501400 524273 502400
rect 495764 499400 496723 501400
rect 498723 499400 499723 501400
rect 501723 499400 502723 501400
rect 504723 499400 505723 501400
rect 507723 499400 508723 501400
rect 510723 499400 511723 501400
rect 513723 499400 514723 501400
rect 516723 499400 517723 501400
rect 519723 500390 524273 501400
rect 528170 500390 528966 510282
rect 519723 499400 528966 500390
rect 495764 498400 528966 499400
rect 495764 496400 496723 498400
rect 498723 496400 499723 498400
rect 501723 496400 502723 498400
rect 504723 496400 505723 498400
rect 507723 496400 508723 498400
rect 510723 496400 511723 498400
rect 513723 496400 514723 498400
rect 516723 496400 517723 498400
rect 519723 496400 528966 498400
rect 495764 495400 528966 496400
rect 495764 493400 496723 495400
rect 498723 493400 499723 495400
rect 501723 493400 502723 495400
rect 504723 493400 505723 495400
rect 507723 493400 508723 495400
rect 510723 493400 511723 495400
rect 513723 493400 514723 495400
rect 516723 493400 517723 495400
rect 519723 493400 528966 495400
rect 495764 492400 528966 493400
rect 495764 490400 496723 492400
rect 498723 490400 499723 492400
rect 501723 490400 502723 492400
rect 504723 490400 505723 492400
rect 507723 490400 508723 492400
rect 510723 490400 511723 492400
rect 513723 490400 514723 492400
rect 516723 490400 517723 492400
rect 519723 490400 528966 492400
rect 495764 489400 528966 490400
rect 495764 487400 496723 489400
rect 498723 487400 499723 489400
rect 501723 487400 502723 489400
rect 504723 487400 505723 489400
rect 507723 487400 508723 489400
rect 510723 487400 511723 489400
rect 513723 487400 514723 489400
rect 516723 487400 517723 489400
rect 519723 487400 528966 489400
rect 495764 486400 528966 487400
rect 43982 483574 44980 486002
rect 495764 484400 496723 486400
rect 498723 484400 499723 486400
rect 501723 484400 502723 486400
rect 504723 484400 505723 486400
rect 507723 484400 508723 486400
rect 510723 484400 511723 486400
rect 513723 484400 514723 486400
rect 516723 484400 517723 486400
rect 519723 484400 528966 486400
rect 43982 483206 46087 483574
rect 43983 483174 46087 483206
rect 495764 483400 528966 484400
rect 43983 482774 45687 483174
rect 495764 481400 496723 483400
rect 498723 481400 499723 483400
rect 501723 481400 502723 483400
rect 504723 481400 505723 483400
rect 507723 481400 508723 483400
rect 510723 481400 511723 483400
rect 513723 481400 514723 483400
rect 516723 481400 517723 483400
rect 519723 481400 528966 483400
rect 495764 480400 528966 481400
rect 495764 478400 496723 480400
rect 498723 478400 499723 480400
rect 501723 478400 502723 480400
rect 504723 478400 505723 480400
rect 507723 478400 508723 480400
rect 510723 478400 511723 480400
rect 513723 478400 514723 480400
rect 516723 478400 517723 480400
rect 519723 478400 528966 480400
rect 495764 477400 528966 478400
rect 495764 475400 496723 477400
rect 498723 475400 499723 477400
rect 501723 475400 502723 477400
rect 504723 475400 505723 477400
rect 507723 475400 508723 477400
rect 510723 475400 511723 477400
rect 513723 475400 514723 477400
rect 516723 475400 517723 477400
rect 519723 475400 528966 477400
rect 495764 474400 528966 475400
rect 495764 472400 496723 474400
rect 498723 472400 499723 474400
rect 501723 472400 502723 474400
rect 504723 472400 505723 474400
rect 507723 472400 508723 474400
rect 510723 472400 511723 474400
rect 513723 472400 514723 474400
rect 516723 472400 517723 474400
rect 519723 472400 528966 474400
rect 495764 471400 528966 472400
rect 495764 469400 496723 471400
rect 498723 469400 499723 471400
rect 501723 469400 502723 471400
rect 504723 469400 505723 471400
rect 507723 469400 508723 471400
rect 510723 469400 511723 471400
rect 513723 469400 514723 471400
rect 516723 469400 517723 471400
rect 519723 469400 528966 471400
rect 495764 468400 528966 469400
rect 495764 466400 496723 468400
rect 498723 466400 499723 468400
rect 501723 466400 502723 468400
rect 504723 466400 505723 468400
rect 507723 466400 508723 468400
rect 510723 466400 511723 468400
rect 513723 466400 514723 468400
rect 516723 466400 517723 468400
rect 519723 466400 528966 468400
rect 495764 465400 528966 466400
rect 495764 463400 496723 465400
rect 498723 463400 499723 465400
rect 501723 463400 502723 465400
rect 504723 463400 505723 465400
rect 507723 463400 508723 465400
rect 510723 463400 511723 465400
rect 513723 463400 514723 465400
rect 516723 463400 517723 465400
rect 519723 463400 528966 465400
rect 495764 462400 528966 463400
rect 495764 460400 496723 462400
rect 498723 460400 499723 462400
rect 501723 460400 502723 462400
rect 504723 460400 505723 462400
rect 507723 460400 508723 462400
rect 510723 460400 511723 462400
rect 513723 460400 514723 462400
rect 516723 460400 517723 462400
rect 519723 460400 528966 462400
rect 495764 459400 528966 460400
rect 495764 457400 496723 459400
rect 498723 457400 499723 459400
rect 501723 457400 502723 459400
rect 504723 457400 505723 459400
rect 507723 457400 508723 459400
rect 510723 457400 511723 459400
rect 513723 457400 514723 459400
rect 516723 457400 517723 459400
rect 519723 457400 528966 459400
rect 495764 456400 528966 457400
rect 495764 454400 496723 456400
rect 498723 454400 499723 456400
rect 501723 454400 502723 456400
rect 504723 454400 505723 456400
rect 507723 454400 508723 456400
rect 510723 454400 511723 456400
rect 513723 454400 514723 456400
rect 516723 454400 517723 456400
rect 519723 454400 528966 456400
rect 495764 453400 528966 454400
rect 495764 451400 496723 453400
rect 498723 451400 499723 453400
rect 501723 451400 502723 453400
rect 504723 451400 505723 453400
rect 507723 451400 508723 453400
rect 510723 451400 511723 453400
rect 513723 451400 514723 453400
rect 516723 451400 517723 453400
rect 519723 451400 528966 453400
rect 495764 450400 528966 451400
rect 495764 448400 496723 450400
rect 498723 448400 499723 450400
rect 501723 448400 502723 450400
rect 504723 448400 505723 450400
rect 507723 448400 508723 450400
rect 510723 448400 511723 450400
rect 513723 448400 514723 450400
rect 516723 448400 517723 450400
rect 519723 448400 528966 450400
rect 495764 447400 528966 448400
rect 495764 445400 496723 447400
rect 498723 445400 499723 447400
rect 501723 445400 502723 447400
rect 504723 445400 505723 447400
rect 507723 445400 508723 447400
rect 510723 445400 511723 447400
rect 513723 445400 514723 447400
rect 516723 445400 517723 447400
rect 519723 445400 528966 447400
rect 495764 444400 528966 445400
rect 495764 442400 496723 444400
rect 498723 442400 499723 444400
rect 501723 442400 502723 444400
rect 504723 442400 505723 444400
rect 507723 442400 508723 444400
rect 510723 442400 511723 444400
rect 513723 442400 514723 444400
rect 516723 442400 517723 444400
rect 519723 442400 528966 444400
rect 495764 441400 528966 442400
rect 495764 439400 496723 441400
rect 498723 439400 499723 441400
rect 501723 439400 502723 441400
rect 504723 439400 505723 441400
rect 507723 439400 508723 441400
rect 510723 439400 511723 441400
rect 513723 439400 514723 441400
rect 516723 439400 517723 441400
rect 519723 439400 528966 441400
rect 495764 438400 528966 439400
rect 495764 436400 496723 438400
rect 498723 436400 499723 438400
rect 501723 436400 502723 438400
rect 504723 436400 505723 438400
rect 507723 436400 508723 438400
rect 510723 436400 511723 438400
rect 513723 436400 514723 438400
rect 516723 436400 517723 438400
rect 519723 436400 528966 438400
rect 495764 435400 528966 436400
rect 495764 433400 496723 435400
rect 498723 433400 499723 435400
rect 501723 433400 502723 435400
rect 504723 433400 505723 435400
rect 507723 433400 508723 435400
rect 510723 433400 511723 435400
rect 513723 433400 514723 435400
rect 516723 433400 517723 435400
rect 519723 433400 528966 435400
rect 495764 422435 528966 433400
rect 402164 377000 495764 378508
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 490208 685800 528967 702351
rect 490208 683800 492200 685800
rect 494200 683800 496200 685800
rect 498200 683800 500200 685800
rect 502200 683800 504200 685800
rect 506200 683800 508200 685800
rect 510200 683800 512200 685800
rect 514200 683800 516200 685800
rect 518200 683800 520200 685800
rect 522200 683800 524200 685800
rect 526200 683800 528967 685800
rect 490208 681800 528967 683800
rect 490208 679800 492200 681800
rect 494200 679800 496200 681800
rect 498200 679800 500200 681800
rect 502200 679800 504200 681800
rect 506200 679800 508200 681800
rect 510200 679800 512200 681800
rect 514200 679800 516200 681800
rect 518200 679800 520200 681800
rect 522200 679800 524200 681800
rect 526200 679800 528967 681800
rect 490208 677800 528967 679800
rect 490208 675800 492200 677800
rect 494200 675800 496200 677800
rect 498200 675800 500200 677800
rect 502200 675800 504200 677800
rect 506200 675800 508200 677800
rect 510200 675800 512200 677800
rect 514200 675800 516200 677800
rect 518200 675800 520200 677800
rect 522200 675800 524200 677800
rect 526200 675800 528967 677800
rect 490208 673800 528967 675800
rect 490208 671800 492200 673800
rect 494200 671800 496200 673800
rect 498200 671800 500200 673800
rect 502200 671800 504200 673800
rect 506200 671800 508200 673800
rect 510200 671800 512200 673800
rect 514200 671800 516200 673800
rect 518200 671800 520200 673800
rect 522200 671800 524200 673800
rect 526200 671800 528967 673800
rect 490208 669800 528967 671800
rect 490208 667800 492200 669800
rect 494200 667800 496200 669800
rect 498200 667800 500200 669800
rect 502200 667800 504200 669800
rect 506200 667800 508200 669800
rect 510200 667800 512200 669800
rect 514200 667800 516200 669800
rect 518200 667800 520200 669800
rect 522200 667800 524200 669800
rect 526200 667800 528967 669800
rect 490208 665800 528967 667800
rect 490208 663800 492200 665800
rect 494200 663800 496200 665800
rect 498200 663800 500200 665800
rect 502200 663800 504200 665800
rect 506200 663800 508200 665800
rect 510200 663800 512200 665800
rect 514200 663800 516200 665800
rect 518200 663800 520200 665800
rect 522200 663800 524200 665800
rect 526200 663800 528967 665800
rect 490208 661800 528967 663800
rect 490208 659800 492200 661800
rect 494200 659800 496200 661800
rect 498200 659800 500200 661800
rect 502200 659800 504200 661800
rect 506200 659800 508200 661800
rect 510200 659800 512200 661800
rect 514200 659800 516200 661800
rect 518200 659800 520200 661800
rect 522200 659800 524200 661800
rect 526200 659800 528967 661800
rect 490208 657800 528967 659800
rect 490208 655800 492200 657800
rect 494200 655800 496200 657800
rect 498200 655800 500200 657800
rect 502200 655800 504200 657800
rect 506200 655800 508200 657800
rect 510200 655800 512200 657800
rect 514200 655800 516200 657800
rect 518200 655800 520200 657800
rect 522200 655800 524200 657800
rect 526200 655800 528967 657800
rect 490208 653800 528967 655800
rect 490208 651800 492200 653800
rect 494200 651800 496200 653800
rect 498200 651800 500200 653800
rect 502200 651800 504200 653800
rect 506200 651800 508200 653800
rect 510200 651800 512200 653800
rect 514200 651800 516200 653800
rect 518200 651800 520200 653800
rect 522200 651800 524200 653800
rect 526200 651800 528967 653800
rect 490208 649800 528967 651800
rect 490208 647800 492200 649800
rect 494200 647800 496200 649800
rect 498200 647800 500200 649800
rect 502200 647800 504200 649800
rect 506200 647800 508200 649800
rect 510200 647800 512200 649800
rect 514200 647800 516200 649800
rect 518200 647800 520200 649800
rect 522200 647800 524200 649800
rect 526200 647800 528967 649800
rect 490208 645800 528967 647800
rect 490208 643800 492200 645800
rect 494200 643800 496200 645800
rect 498200 643800 500200 645800
rect 502200 643800 504200 645800
rect 506200 643800 508200 645800
rect 510200 643800 512200 645800
rect 514200 643800 516200 645800
rect 518200 643800 520200 645800
rect 522200 643800 524200 645800
rect 526200 643800 528967 645800
rect 490208 641800 528967 643800
rect 490208 639800 492200 641800
rect 494200 639800 496200 641800
rect 498200 639800 500200 641800
rect 502200 639800 504200 641800
rect 506200 639800 508200 641800
rect 510200 639800 512200 641800
rect 514200 639800 516200 641800
rect 518200 639800 520200 641800
rect 522200 639800 524200 641800
rect 526200 639800 528967 641800
rect 490208 637800 528967 639800
rect 490208 635800 492200 637800
rect 494200 635800 496200 637800
rect 498200 635800 500200 637800
rect 502200 635800 504200 637800
rect 506200 635800 508200 637800
rect 510200 635800 512200 637800
rect 514200 635800 516200 637800
rect 518200 635800 520200 637800
rect 522200 635800 524200 637800
rect 526200 635800 528967 637800
rect 490208 633800 528967 635800
rect 490208 631800 492200 633800
rect 494200 631800 496200 633800
rect 498200 631800 500200 633800
rect 502200 631800 504200 633800
rect 506200 631800 508200 633800
rect 510200 631800 512200 633800
rect 514200 631800 516200 633800
rect 518200 631800 520200 633800
rect 522200 631800 524200 633800
rect 526200 631800 528967 633800
rect 326401 630473 327081 631055
rect 490208 629800 528967 631800
rect 490208 627800 492200 629800
rect 494200 627800 496200 629800
rect 498200 627800 500200 629800
rect 502200 627800 504200 629800
rect 506200 627800 508200 629800
rect 510200 627800 512200 629800
rect 514200 627800 516200 629800
rect 518200 627800 520200 629800
rect 522200 627800 524200 629800
rect 526200 627800 528967 629800
rect 490208 625800 528967 627800
rect 490208 623800 492200 625800
rect 494200 623800 496200 625800
rect 498200 623800 500200 625800
rect 502200 623800 504200 625800
rect 506200 623800 508200 625800
rect 510200 623800 512200 625800
rect 514200 623800 516200 625800
rect 518200 623800 520200 625800
rect 522200 623800 524200 625800
rect 526200 623800 528967 625800
rect 490208 621800 528967 623800
rect 490208 619800 492200 621800
rect 494200 619800 496200 621800
rect 498200 619800 500200 621800
rect 502200 619800 504200 621800
rect 506200 619800 508200 621800
rect 510200 619800 512200 621800
rect 514200 619800 516200 621800
rect 518200 619800 520200 621800
rect 522200 619800 524200 621800
rect 526200 619800 528967 621800
rect 490208 617800 528967 619800
rect 490208 615800 492200 617800
rect 494200 615800 496200 617800
rect 498200 615800 500200 617800
rect 502200 615800 504200 617800
rect 506200 615800 508200 617800
rect 510200 615800 512200 617800
rect 514200 615800 516200 617800
rect 518200 615800 520200 617800
rect 522200 615800 524200 617800
rect 526200 615800 528967 617800
rect 490208 613800 528967 615800
rect 490208 611800 492200 613800
rect 494200 611800 496200 613800
rect 498200 611800 500200 613800
rect 502200 611800 504200 613800
rect 506200 611800 508200 613800
rect 510200 611800 512200 613800
rect 514200 611800 516200 613800
rect 518200 611800 520200 613800
rect 522200 611800 524200 613800
rect 526200 611800 528967 613800
rect 490208 609800 528967 611800
rect 490208 607800 492200 609800
rect 494200 607800 496200 609800
rect 498200 607800 500200 609800
rect 502200 607800 504200 609800
rect 506200 607800 508200 609800
rect 510200 607800 512200 609800
rect 514200 607800 516200 609800
rect 518200 607800 520200 609800
rect 522200 607800 524200 609800
rect 526200 607800 528967 609800
rect 490208 605800 528967 607800
rect 490208 603800 492200 605800
rect 494200 603800 496200 605800
rect 498200 603800 500200 605800
rect 502200 603800 504200 605800
rect 506200 603800 508200 605800
rect 510200 603800 512200 605800
rect 514200 603800 516200 605800
rect 518200 603800 520200 605800
rect 522200 603800 524200 605800
rect 526200 603800 528967 605800
rect 490208 601800 528967 603800
rect 490208 599800 492200 601800
rect 494200 599800 496200 601800
rect 498200 599800 500200 601800
rect 502200 599800 504200 601800
rect 506200 599800 508200 601800
rect 510200 599800 512200 601800
rect 514200 599800 516200 601800
rect 518200 599800 520200 601800
rect 522200 599800 524200 601800
rect 526200 599800 528967 601800
rect 490208 597800 528967 599800
rect 490208 595800 492200 597800
rect 494200 595800 496200 597800
rect 498200 595800 500200 597800
rect 502200 595800 504200 597800
rect 506200 595800 508200 597800
rect 510200 595800 512200 597800
rect 514200 595800 516200 597800
rect 518200 595800 520200 597800
rect 522200 595800 524200 597800
rect 526200 595800 528967 597800
rect 490208 593800 528967 595800
rect 490208 591800 492200 593800
rect 494200 591800 496200 593800
rect 498200 591800 500200 593800
rect 502200 591800 504200 593800
rect 506200 591800 508200 593800
rect 510200 591800 512200 593800
rect 514200 591800 516200 593800
rect 518200 591800 520200 593800
rect 522200 591800 524200 593800
rect 526200 591800 528967 593800
rect 490208 589800 528967 591800
rect 490208 587800 492200 589800
rect 494200 587800 496200 589800
rect 498200 587800 500200 589800
rect 502200 587800 504200 589800
rect 506200 587800 508200 589800
rect 510200 587800 512200 589800
rect 514200 587800 516200 589800
rect 518200 587800 520200 589800
rect 522200 587800 524200 589800
rect 526200 587800 528967 589800
rect 203279 565294 215403 581258
rect 490208 551657 528967 587800
rect 490208 549657 491621 551657
rect 493621 549657 494621 551657
rect 496621 549657 497621 551657
rect 499621 549657 500621 551657
rect 502621 549657 503621 551657
rect 505621 549657 506621 551657
rect 508621 549657 509621 551657
rect 511621 549657 512621 551657
rect 514621 549657 515621 551657
rect 517621 549657 518621 551657
rect 520621 549657 528967 551657
rect 490208 548657 528967 549657
rect 490208 546657 491621 548657
rect 493621 546657 494621 548657
rect 496621 546657 497621 548657
rect 499621 546657 500621 548657
rect 502621 546657 503621 548657
rect 505621 546657 506621 548657
rect 508621 546657 509621 548657
rect 511621 546657 512621 548657
rect 514621 546657 515621 548657
rect 517621 546657 518621 548657
rect 520621 546657 528967 548657
rect 490208 545657 528967 546657
rect 490208 543657 491621 545657
rect 493621 543657 494621 545657
rect 496621 543657 497621 545657
rect 499621 543657 500621 545657
rect 502621 543657 503621 545657
rect 505621 543657 506621 545657
rect 508621 543657 509621 545657
rect 511621 543657 512621 545657
rect 514621 543657 515621 545657
rect 517621 543657 518621 545657
rect 520621 543657 528967 545657
rect 490208 542657 528967 543657
rect 490208 540657 491621 542657
rect 493621 540657 494621 542657
rect 496621 540657 497621 542657
rect 499621 540657 500621 542657
rect 502621 540657 503621 542657
rect 505621 540657 506621 542657
rect 508621 540657 509621 542657
rect 511621 540657 512621 542657
rect 514621 540657 515621 542657
rect 517621 540657 518621 542657
rect 520621 540657 528967 542657
rect 490208 539657 528967 540657
rect 490208 537657 491621 539657
rect 493621 537657 494621 539657
rect 496621 537657 497621 539657
rect 499621 537657 500621 539657
rect 502621 537657 503621 539657
rect 505621 537657 506621 539657
rect 508621 537657 509621 539657
rect 511621 537657 512621 539657
rect 514621 537657 515621 539657
rect 517621 537657 518621 539657
rect 520621 537657 528967 539657
rect 490208 536657 528967 537657
rect 490208 534657 491621 536657
rect 493621 534657 494621 536657
rect 496621 534657 497621 536657
rect 499621 534657 500621 536657
rect 502621 534657 503621 536657
rect 505621 534657 506621 536657
rect 508621 534657 509621 536657
rect 511621 534657 512621 536657
rect 514621 534657 515621 536657
rect 517621 534657 518621 536657
rect 520621 534657 528967 536657
rect 490208 533657 528967 534657
rect 490208 531657 491621 533657
rect 493621 531657 494621 533657
rect 496621 531657 497621 533657
rect 499621 531657 500621 533657
rect 502621 531657 503621 533657
rect 505621 531657 506621 533657
rect 508621 531657 509621 533657
rect 511621 531657 512621 533657
rect 514621 531657 515621 533657
rect 517621 531657 518621 533657
rect 520621 531657 528967 533657
rect 490208 530657 528967 531657
rect 490208 528657 491621 530657
rect 493621 528657 494621 530657
rect 496621 528657 497621 530657
rect 499621 528657 500621 530657
rect 502621 528657 503621 530657
rect 505621 528657 506621 530657
rect 508621 528657 509621 530657
rect 511621 528657 512621 530657
rect 514621 528657 515621 530657
rect 517621 528657 518621 530657
rect 520621 528657 528967 530657
rect 490208 527657 528967 528657
rect 490208 527108 491621 527657
rect 493621 527108 494621 527657
rect 402164 525657 495764 527108
rect 496621 525657 497621 527657
rect 499621 525657 500621 527657
rect 502621 525657 503621 527657
rect 505621 525657 506621 527657
rect 508621 525657 509621 527657
rect 511621 525657 512621 527657
rect 514621 525657 515621 527657
rect 517621 525657 518621 527657
rect 520621 525657 528967 527657
rect 402164 524657 528967 525657
rect 402164 522657 495764 524657
rect 496621 522657 497621 524657
rect 499621 522657 500621 524657
rect 502621 522657 503621 524657
rect 505621 522657 506621 524657
rect 508621 522657 509621 524657
rect 511621 522657 512621 524657
rect 514621 522657 515621 524657
rect 517621 522657 518621 524657
rect 520621 522657 528967 524657
rect 402164 521657 528967 522657
rect 402164 521462 495764 521657
rect 402164 519462 421473 521462
rect 423473 519462 424473 521462
rect 426473 519462 427473 521462
rect 429473 519462 430473 521462
rect 432473 519462 433473 521462
rect 435473 519462 436473 521462
rect 438473 519462 439473 521462
rect 441473 519462 442473 521462
rect 444473 519462 445473 521462
rect 447473 519462 448473 521462
rect 450473 519462 451473 521462
rect 453473 519462 454473 521462
rect 456473 519462 457473 521462
rect 459473 519462 460473 521462
rect 462473 519462 463473 521462
rect 465473 519462 466473 521462
rect 468473 519462 469473 521462
rect 471473 519462 472473 521462
rect 474473 519657 495764 521462
rect 496621 519657 497621 521657
rect 499621 519657 500621 521657
rect 502621 519657 503621 521657
rect 505621 519657 506621 521657
rect 508621 519657 509621 521657
rect 511621 519657 512621 521657
rect 514621 519657 515621 521657
rect 517621 519657 518621 521657
rect 520621 519657 528967 521657
rect 474473 519462 528967 519657
rect 402164 518657 528967 519462
rect 402164 518462 495764 518657
rect 402164 516462 421473 518462
rect 423473 516462 424473 518462
rect 426473 516462 427473 518462
rect 429473 516462 430473 518462
rect 432473 516462 433473 518462
rect 435473 516462 436473 518462
rect 438473 516462 439473 518462
rect 441473 516462 442473 518462
rect 444473 516462 445473 518462
rect 447473 516462 448473 518462
rect 450473 516462 451473 518462
rect 453473 516462 454473 518462
rect 456473 516462 457473 518462
rect 459473 516462 460473 518462
rect 462473 516462 463473 518462
rect 465473 516462 466473 518462
rect 468473 516462 469473 518462
rect 471473 516462 472473 518462
rect 474473 516657 495764 518462
rect 496621 516657 497621 518657
rect 499621 516657 500621 518657
rect 502621 516657 503621 518657
rect 505621 516657 506621 518657
rect 508621 516657 509621 518657
rect 511621 516657 512621 518657
rect 514621 516657 515621 518657
rect 517621 516657 518621 518657
rect 520621 516657 528967 518657
rect 474473 516462 528967 516657
rect 402164 515657 528967 516462
rect 402164 515462 495764 515657
rect 402164 513462 421473 515462
rect 423473 513462 424473 515462
rect 426473 513462 427473 515462
rect 429473 513462 430473 515462
rect 432473 513462 433473 515462
rect 435473 513462 436473 515462
rect 438473 513462 439473 515462
rect 441473 513462 442473 515462
rect 444473 513462 445473 515462
rect 447473 513462 448473 515462
rect 450473 513462 451473 515462
rect 453473 513462 454473 515462
rect 456473 513462 457473 515462
rect 459473 513462 460473 515462
rect 462473 513462 463473 515462
rect 465473 513462 466473 515462
rect 468473 513462 469473 515462
rect 471473 513462 472473 515462
rect 474473 513657 495764 515462
rect 496621 513657 497621 515657
rect 499621 513657 500621 515657
rect 502621 513657 503621 515657
rect 505621 513657 506621 515657
rect 508621 513657 509621 515657
rect 511621 513657 512621 515657
rect 514621 513657 515621 515657
rect 517621 513657 518621 515657
rect 520621 513657 528967 515657
rect 474473 513462 528967 513657
rect 402164 512657 528967 513462
rect 402164 512462 495764 512657
rect 402164 510462 421473 512462
rect 423473 510462 424473 512462
rect 426473 510462 427473 512462
rect 429473 510462 430473 512462
rect 432473 510462 433473 512462
rect 435473 510462 436473 512462
rect 438473 510462 439473 512462
rect 441473 510462 442473 512462
rect 444473 510462 445473 512462
rect 447473 510462 448473 512462
rect 450473 510462 451473 512462
rect 453473 510462 454473 512462
rect 456473 510462 457473 512462
rect 459473 510462 460473 512462
rect 462473 510462 463473 512462
rect 465473 510462 466473 512462
rect 468473 510462 469473 512462
rect 471473 510462 472473 512462
rect 474473 510657 495764 512462
rect 496621 510657 497621 512657
rect 499621 510657 500621 512657
rect 502621 510657 503621 512657
rect 505621 510657 506621 512657
rect 508621 510657 509621 512657
rect 511621 510657 512621 512657
rect 514621 510657 515621 512657
rect 517621 510657 518621 512657
rect 520621 510657 528967 512657
rect 474473 510462 528967 510657
rect 402164 509657 528967 510462
rect 402164 509462 495764 509657
rect 402164 507462 421473 509462
rect 423473 507462 424473 509462
rect 426473 507462 427473 509462
rect 429473 507462 430473 509462
rect 432473 507462 433473 509462
rect 435473 507462 436473 509462
rect 438473 507462 439473 509462
rect 441473 507462 442473 509462
rect 444473 507462 445473 509462
rect 447473 507462 448473 509462
rect 450473 507462 451473 509462
rect 453473 507462 454473 509462
rect 456473 507462 457473 509462
rect 459473 507462 460473 509462
rect 462473 507462 463473 509462
rect 465473 507462 466473 509462
rect 468473 507462 469473 509462
rect 471473 507462 472473 509462
rect 474473 507657 495764 509462
rect 496621 507657 497621 509657
rect 499621 507657 500621 509657
rect 502621 507657 503621 509657
rect 505621 507657 506621 509657
rect 508621 507657 509621 509657
rect 511621 507657 512621 509657
rect 514621 507657 515621 509657
rect 517621 507657 518621 509657
rect 520621 507657 528967 509657
rect 474473 507462 528967 507657
rect 402164 506657 528967 507462
rect 402164 506462 495764 506657
rect 402164 504462 421473 506462
rect 423473 504462 424473 506462
rect 426473 504462 427473 506462
rect 429473 504462 430473 506462
rect 432473 504462 433473 506462
rect 435473 504462 436473 506462
rect 438473 504462 439473 506462
rect 441473 504462 442473 506462
rect 444473 504462 445473 506462
rect 447473 504462 448473 506462
rect 450473 504462 451473 506462
rect 453473 504462 454473 506462
rect 456473 504462 457473 506462
rect 459473 504462 460473 506462
rect 462473 504462 463473 506462
rect 465473 504462 466473 506462
rect 468473 504462 469473 506462
rect 471473 504462 472473 506462
rect 474473 504657 495764 506462
rect 496621 504657 497621 506657
rect 499621 504657 500621 506657
rect 502621 504657 503621 506657
rect 505621 504657 506621 506657
rect 508621 504657 509621 506657
rect 511621 504657 512621 506657
rect 514621 504657 515621 506657
rect 517621 504657 518621 506657
rect 520621 504657 528967 506657
rect 474473 504462 528967 504657
rect 402164 503657 528967 504462
rect 402164 503462 495764 503657
rect 402164 501462 421473 503462
rect 423473 501462 424473 503462
rect 426473 501462 427473 503462
rect 429473 501462 430473 503462
rect 432473 501462 433473 503462
rect 435473 501462 436473 503462
rect 438473 501462 439473 503462
rect 441473 501462 442473 503462
rect 444473 501462 445473 503462
rect 447473 501462 448473 503462
rect 450473 501462 451473 503462
rect 453473 501462 454473 503462
rect 456473 501462 457473 503462
rect 459473 501462 460473 503462
rect 462473 501462 463473 503462
rect 465473 501462 466473 503462
rect 468473 501462 469473 503462
rect 471473 501462 472473 503462
rect 474473 501657 495764 503462
rect 496621 501657 497621 503657
rect 499621 501657 500621 503657
rect 502621 501657 503621 503657
rect 505621 501657 506621 503657
rect 508621 501657 509621 503657
rect 511621 501657 512621 503657
rect 514621 501657 515621 503657
rect 517621 501657 518621 503657
rect 520621 501657 528967 503657
rect 474473 501462 528967 501657
rect 402164 500657 528967 501462
rect 402164 500462 495764 500657
rect 402164 498462 421473 500462
rect 423473 498462 424473 500462
rect 426473 498462 427473 500462
rect 429473 498462 430473 500462
rect 432473 498462 433473 500462
rect 435473 498462 436473 500462
rect 438473 498462 439473 500462
rect 441473 498462 442473 500462
rect 444473 498462 445473 500462
rect 447473 498462 448473 500462
rect 450473 498462 451473 500462
rect 453473 498462 454473 500462
rect 456473 498462 457473 500462
rect 459473 498462 460473 500462
rect 462473 498462 463473 500462
rect 465473 498462 466473 500462
rect 468473 498462 469473 500462
rect 471473 498462 472473 500462
rect 474473 498657 495764 500462
rect 496621 498657 497621 500657
rect 499621 498657 500621 500657
rect 502621 498657 503621 500657
rect 505621 498657 506621 500657
rect 508621 498657 509621 500657
rect 511621 498657 512621 500657
rect 514621 498657 515621 500657
rect 517621 498657 518621 500657
rect 520621 498657 528967 500657
rect 474473 498462 528967 498657
rect 402164 497657 528967 498462
rect 402164 497462 495764 497657
rect 402164 495462 421473 497462
rect 423473 495462 424473 497462
rect 426473 495462 427473 497462
rect 429473 495462 430473 497462
rect 432473 495462 433473 497462
rect 435473 495462 436473 497462
rect 438473 495462 439473 497462
rect 441473 495462 442473 497462
rect 444473 495462 445473 497462
rect 447473 495462 448473 497462
rect 450473 495462 451473 497462
rect 453473 495462 454473 497462
rect 456473 495462 457473 497462
rect 459473 495462 460473 497462
rect 462473 495462 463473 497462
rect 465473 495462 466473 497462
rect 468473 495462 469473 497462
rect 471473 495462 472473 497462
rect 474473 495657 495764 497462
rect 496621 495657 497621 497657
rect 499621 495657 500621 497657
rect 502621 495657 503621 497657
rect 505621 495657 506621 497657
rect 508621 495657 509621 497657
rect 511621 495657 512621 497657
rect 514621 495657 515621 497657
rect 517621 495657 518621 497657
rect 520621 495657 528967 497657
rect 474473 495462 528967 495657
rect 402164 494657 528967 495462
rect 402164 494462 495764 494657
rect 402164 492462 421473 494462
rect 423473 492462 424473 494462
rect 426473 492462 427473 494462
rect 429473 492462 430473 494462
rect 432473 492462 433473 494462
rect 435473 492462 436473 494462
rect 438473 492462 439473 494462
rect 441473 492462 442473 494462
rect 444473 492462 445473 494462
rect 447473 492462 448473 494462
rect 450473 492462 451473 494462
rect 453473 492462 454473 494462
rect 456473 492462 457473 494462
rect 459473 492462 460473 494462
rect 462473 492462 463473 494462
rect 465473 492462 466473 494462
rect 468473 492462 469473 494462
rect 471473 492462 472473 494462
rect 474473 492657 495764 494462
rect 496621 492657 497621 494657
rect 499621 492657 500621 494657
rect 502621 492657 503621 494657
rect 505621 492657 506621 494657
rect 508621 492657 509621 494657
rect 511621 492657 512621 494657
rect 514621 492657 515621 494657
rect 517621 492657 518621 494657
rect 520621 492657 528967 494657
rect 474473 492462 528967 492657
rect 402164 491657 528967 492462
rect 402164 491462 495764 491657
rect 402164 489462 421473 491462
rect 423473 489462 424473 491462
rect 426473 489462 427473 491462
rect 429473 489462 430473 491462
rect 432473 489462 433473 491462
rect 435473 489462 436473 491462
rect 438473 489462 439473 491462
rect 441473 489462 442473 491462
rect 444473 489462 445473 491462
rect 447473 489462 448473 491462
rect 450473 489462 451473 491462
rect 453473 489462 454473 491462
rect 456473 489462 457473 491462
rect 459473 489462 460473 491462
rect 462473 489462 463473 491462
rect 465473 489462 466473 491462
rect 468473 489462 469473 491462
rect 471473 489462 472473 491462
rect 474473 489657 495764 491462
rect 496621 489657 497621 491657
rect 499621 489657 500621 491657
rect 502621 489657 503621 491657
rect 505621 489657 506621 491657
rect 508621 489657 509621 491657
rect 511621 489657 512621 491657
rect 514621 489657 515621 491657
rect 517621 489657 518621 491657
rect 520621 489657 528967 491657
rect 474473 489462 528967 489657
rect 402164 488657 528967 489462
rect 402164 488462 495764 488657
rect 402164 486462 421473 488462
rect 423473 486462 424473 488462
rect 426473 486462 427473 488462
rect 429473 486462 430473 488462
rect 432473 486462 433473 488462
rect 435473 486462 436473 488462
rect 438473 486462 439473 488462
rect 441473 486462 442473 488462
rect 444473 486462 445473 488462
rect 447473 486462 448473 488462
rect 450473 486462 451473 488462
rect 453473 486462 454473 488462
rect 456473 486462 457473 488462
rect 459473 486462 460473 488462
rect 462473 486462 463473 488462
rect 465473 486462 466473 488462
rect 468473 486462 469473 488462
rect 471473 486462 472473 488462
rect 474473 486657 495764 488462
rect 496621 486657 497621 488657
rect 499621 486657 500621 488657
rect 502621 486657 503621 488657
rect 505621 486657 506621 488657
rect 508621 486657 509621 488657
rect 511621 486657 512621 488657
rect 514621 486657 515621 488657
rect 517621 486657 518621 488657
rect 520621 486657 528967 488657
rect 474473 486462 528967 486657
rect 402164 485657 528967 486462
rect 402164 485462 495764 485657
rect 402164 483462 421473 485462
rect 423473 483462 424473 485462
rect 426473 483462 427473 485462
rect 429473 483462 430473 485462
rect 432473 483462 433473 485462
rect 435473 483462 436473 485462
rect 438473 483462 439473 485462
rect 441473 483462 442473 485462
rect 444473 483462 445473 485462
rect 447473 483462 448473 485462
rect 450473 483462 451473 485462
rect 453473 483462 454473 485462
rect 456473 483462 457473 485462
rect 459473 483462 460473 485462
rect 462473 483462 463473 485462
rect 465473 483462 466473 485462
rect 468473 483462 469473 485462
rect 471473 483462 472473 485462
rect 474473 483657 495764 485462
rect 496621 483657 497621 485657
rect 499621 483657 500621 485657
rect 502621 483657 503621 485657
rect 505621 483657 506621 485657
rect 508621 483657 509621 485657
rect 511621 483657 512621 485657
rect 514621 483657 515621 485657
rect 517621 483657 518621 485657
rect 520621 483657 528967 485657
rect 474473 483462 528967 483657
rect 402164 482657 528967 483462
rect 402164 482462 495764 482657
rect 402164 480462 421473 482462
rect 423473 480462 424473 482462
rect 426473 480462 427473 482462
rect 429473 480462 430473 482462
rect 432473 480462 433473 482462
rect 435473 480462 436473 482462
rect 438473 480462 439473 482462
rect 441473 480462 442473 482462
rect 444473 480462 445473 482462
rect 447473 480462 448473 482462
rect 450473 480462 451473 482462
rect 453473 480462 454473 482462
rect 456473 480462 457473 482462
rect 459473 480462 460473 482462
rect 462473 480462 463473 482462
rect 465473 480462 466473 482462
rect 468473 480462 469473 482462
rect 471473 480462 472473 482462
rect 474473 480657 495764 482462
rect 496621 480657 497621 482657
rect 499621 480657 500621 482657
rect 502621 480657 503621 482657
rect 505621 480657 506621 482657
rect 508621 480657 509621 482657
rect 511621 480657 512621 482657
rect 514621 480657 515621 482657
rect 517621 480657 518621 482657
rect 520621 480657 528967 482657
rect 474473 480462 528967 480657
rect 402164 479657 528967 480462
rect 402164 479462 495764 479657
rect 402164 477462 421473 479462
rect 423473 477462 424473 479462
rect 426473 477462 427473 479462
rect 429473 477462 430473 479462
rect 432473 477462 433473 479462
rect 435473 477462 436473 479462
rect 438473 477462 439473 479462
rect 441473 477462 442473 479462
rect 444473 477462 445473 479462
rect 447473 477462 448473 479462
rect 450473 477462 451473 479462
rect 453473 477462 454473 479462
rect 456473 477462 457473 479462
rect 459473 477462 460473 479462
rect 462473 477462 463473 479462
rect 465473 477462 466473 479462
rect 468473 477462 469473 479462
rect 471473 477462 472473 479462
rect 474473 477657 495764 479462
rect 496621 477657 497621 479657
rect 499621 477657 500621 479657
rect 502621 477657 503621 479657
rect 505621 477657 506621 479657
rect 508621 477657 509621 479657
rect 511621 477657 512621 479657
rect 514621 477657 515621 479657
rect 517621 477657 518621 479657
rect 520621 477657 528967 479657
rect 474473 477462 528967 477657
rect 402164 476657 528967 477462
rect 402164 476462 495764 476657
rect 402164 474462 421473 476462
rect 423473 474462 424473 476462
rect 426473 474462 427473 476462
rect 429473 474462 430473 476462
rect 432473 474462 433473 476462
rect 435473 474462 436473 476462
rect 438473 474462 439473 476462
rect 441473 474462 442473 476462
rect 444473 474462 445473 476462
rect 447473 474462 448473 476462
rect 450473 474462 451473 476462
rect 453473 474462 454473 476462
rect 456473 474462 457473 476462
rect 459473 474462 460473 476462
rect 462473 474462 463473 476462
rect 465473 474462 466473 476462
rect 468473 474462 469473 476462
rect 471473 474462 472473 476462
rect 474473 474657 495764 476462
rect 496621 474657 497621 476657
rect 499621 474657 500621 476657
rect 502621 474657 503621 476657
rect 505621 474657 506621 476657
rect 508621 474657 509621 476657
rect 511621 474657 512621 476657
rect 514621 474657 515621 476657
rect 517621 474657 518621 476657
rect 520621 474657 528967 476657
rect 474473 474462 528967 474657
rect 402164 473657 528967 474462
rect 402164 473462 495764 473657
rect 402164 471462 421473 473462
rect 423473 471462 424473 473462
rect 426473 471462 427473 473462
rect 429473 471462 430473 473462
rect 432473 471462 433473 473462
rect 435473 471462 436473 473462
rect 438473 471462 439473 473462
rect 441473 471462 442473 473462
rect 444473 471462 445473 473462
rect 447473 471462 448473 473462
rect 450473 471462 451473 473462
rect 453473 471462 454473 473462
rect 456473 471462 457473 473462
rect 459473 471462 460473 473462
rect 462473 471462 463473 473462
rect 465473 471462 466473 473462
rect 468473 471462 469473 473462
rect 471473 471462 472473 473462
rect 474473 471657 495764 473462
rect 496621 471657 497621 473657
rect 499621 471657 500621 473657
rect 502621 471657 503621 473657
rect 505621 471657 506621 473657
rect 508621 471657 509621 473657
rect 511621 471657 512621 473657
rect 514621 471657 515621 473657
rect 517621 471657 518621 473657
rect 520621 471657 528967 473657
rect 474473 471462 528967 471657
rect 402164 470657 528967 471462
rect 402164 470462 495764 470657
rect 402164 468462 421473 470462
rect 423473 468462 424473 470462
rect 426473 468462 427473 470462
rect 429473 468462 430473 470462
rect 432473 468462 433473 470462
rect 435473 468462 436473 470462
rect 438473 468462 439473 470462
rect 441473 468462 442473 470462
rect 444473 468462 445473 470462
rect 447473 468462 448473 470462
rect 450473 468462 451473 470462
rect 453473 468462 454473 470462
rect 456473 468462 457473 470462
rect 459473 468462 460473 470462
rect 462473 468462 463473 470462
rect 465473 468462 466473 470462
rect 468473 468462 469473 470462
rect 471473 468462 472473 470462
rect 474473 468657 495764 470462
rect 496621 468657 497621 470657
rect 499621 468657 500621 470657
rect 502621 468657 503621 470657
rect 505621 468657 506621 470657
rect 508621 468657 509621 470657
rect 511621 468657 512621 470657
rect 514621 468657 515621 470657
rect 517621 468657 518621 470657
rect 520621 468657 528967 470657
rect 474473 468462 528967 468657
rect 402164 467657 528967 468462
rect 402164 467462 495764 467657
rect 402164 465462 421473 467462
rect 423473 465462 424473 467462
rect 426473 465462 427473 467462
rect 429473 465462 430473 467462
rect 432473 465462 433473 467462
rect 435473 465462 436473 467462
rect 438473 465462 439473 467462
rect 441473 465462 442473 467462
rect 444473 465462 445473 467462
rect 447473 465462 448473 467462
rect 450473 465462 451473 467462
rect 453473 465462 454473 467462
rect 456473 465462 457473 467462
rect 459473 465462 460473 467462
rect 462473 465462 463473 467462
rect 465473 465462 466473 467462
rect 468473 465462 469473 467462
rect 471473 465462 472473 467462
rect 474473 465657 495764 467462
rect 496621 465657 497621 467657
rect 499621 465657 500621 467657
rect 502621 465657 503621 467657
rect 505621 465657 506621 467657
rect 508621 465657 509621 467657
rect 511621 465657 512621 467657
rect 514621 465657 515621 467657
rect 517621 465657 518621 467657
rect 520621 465657 528967 467657
rect 474473 465462 528967 465657
rect 402164 464657 528967 465462
rect 402164 464462 495764 464657
rect 402164 462462 421473 464462
rect 423473 462462 424473 464462
rect 426473 462462 427473 464462
rect 429473 462462 430473 464462
rect 432473 462462 433473 464462
rect 435473 462462 436473 464462
rect 438473 462462 439473 464462
rect 441473 462462 442473 464462
rect 444473 462462 445473 464462
rect 447473 462462 448473 464462
rect 450473 462462 451473 464462
rect 453473 462462 454473 464462
rect 456473 462462 457473 464462
rect 459473 462462 460473 464462
rect 462473 462462 463473 464462
rect 465473 462462 466473 464462
rect 468473 462462 469473 464462
rect 471473 462462 472473 464462
rect 474473 462657 495764 464462
rect 496621 462657 497621 464657
rect 499621 462657 500621 464657
rect 502621 462657 503621 464657
rect 505621 462657 506621 464657
rect 508621 462657 509621 464657
rect 511621 462657 512621 464657
rect 514621 462657 515621 464657
rect 517621 462657 518621 464657
rect 520621 462657 528967 464657
rect 474473 462462 528967 462657
rect 402164 461657 528967 462462
rect 402164 461462 495764 461657
rect 402164 459462 421473 461462
rect 423473 459462 424473 461462
rect 426473 459462 427473 461462
rect 429473 459462 430473 461462
rect 432473 459462 433473 461462
rect 435473 459462 436473 461462
rect 438473 459462 439473 461462
rect 441473 459462 442473 461462
rect 444473 459462 445473 461462
rect 447473 459462 448473 461462
rect 450473 459462 451473 461462
rect 453473 459462 454473 461462
rect 456473 459462 457473 461462
rect 459473 459462 460473 461462
rect 462473 459462 463473 461462
rect 465473 459462 466473 461462
rect 468473 459462 469473 461462
rect 471473 459462 472473 461462
rect 474473 459657 495764 461462
rect 496621 459657 497621 461657
rect 499621 459657 500621 461657
rect 502621 459657 503621 461657
rect 505621 459657 506621 461657
rect 508621 459657 509621 461657
rect 511621 459657 512621 461657
rect 514621 459657 515621 461657
rect 517621 459657 518621 461657
rect 520621 459657 528967 461657
rect 474473 459462 528967 459657
rect 402164 458657 528967 459462
rect 402164 458462 495764 458657
rect 402164 456462 421473 458462
rect 423473 456462 424473 458462
rect 426473 456462 427473 458462
rect 429473 456462 430473 458462
rect 432473 456462 433473 458462
rect 435473 456462 436473 458462
rect 438473 456462 439473 458462
rect 441473 456462 442473 458462
rect 444473 456462 445473 458462
rect 447473 456462 448473 458462
rect 450473 456462 451473 458462
rect 453473 456462 454473 458462
rect 456473 456462 457473 458462
rect 459473 456462 460473 458462
rect 462473 456462 463473 458462
rect 465473 456462 466473 458462
rect 468473 456462 469473 458462
rect 471473 456462 472473 458462
rect 474473 456657 495764 458462
rect 496621 456657 497621 458657
rect 499621 456657 500621 458657
rect 502621 456657 503621 458657
rect 505621 456657 506621 458657
rect 508621 456657 509621 458657
rect 511621 456657 512621 458657
rect 514621 456657 515621 458657
rect 517621 456657 518621 458657
rect 520621 456657 528967 458657
rect 474473 456462 528967 456657
rect 402164 455657 528967 456462
rect 402164 453657 495764 455657
rect 496621 453657 497621 455657
rect 499621 453657 500621 455657
rect 502621 453657 503621 455657
rect 505621 453657 506621 455657
rect 508621 453657 509621 455657
rect 511621 453657 512621 455657
rect 514621 453657 515621 455657
rect 517621 453657 518621 455657
rect 520621 453657 528967 455657
rect 402164 452657 528967 453657
rect 402164 450657 495764 452657
rect 496621 450657 497621 452657
rect 499621 450657 500621 452657
rect 502621 450657 503621 452657
rect 505621 450657 506621 452657
rect 508621 450657 509621 452657
rect 511621 450657 512621 452657
rect 514621 450657 515621 452657
rect 517621 450657 518621 452657
rect 520621 450657 528967 452657
rect 402164 449657 528967 450657
rect 402164 447657 495764 449657
rect 496621 447657 497621 449657
rect 499621 447657 500621 449657
rect 502621 447657 503621 449657
rect 505621 447657 506621 449657
rect 508621 447657 509621 449657
rect 511621 447657 512621 449657
rect 514621 447657 515621 449657
rect 517621 447657 518621 449657
rect 520621 447657 528967 449657
rect 402164 446657 528967 447657
rect 402164 444657 495764 446657
rect 496621 444657 497621 446657
rect 499621 444657 500621 446657
rect 502621 444657 503621 446657
rect 505621 444657 506621 446657
rect 508621 444657 509621 446657
rect 511621 444657 512621 446657
rect 514621 444657 515621 446657
rect 517621 444657 518621 446657
rect 520621 444657 528967 446657
rect 402164 443657 528967 444657
rect 402164 441657 495764 443657
rect 496621 441657 497621 443657
rect 499621 441657 500621 443657
rect 502621 441657 503621 443657
rect 505621 441657 506621 443657
rect 508621 441657 509621 443657
rect 511621 441657 512621 443657
rect 514621 441657 515621 443657
rect 517621 441657 518621 443657
rect 520621 441657 528967 443657
rect 402164 422443 528967 441657
rect 402164 419444 495764 422443
use Cascode_Amp  Cascode_Amp_0
timestamp 1669601918
transform 0 -1 166000 1 0 311422
box -28448 -26417 68466 42615
use Cascode_Amp  Cascode_Amp_1
timestamp 1669601918
transform 0 -1 166000 1 0 448972
box -28448 -26417 68466 42615
use LNA_final  LNA_final_0
timestamp 1669601918
transform 0 1 404562 -1 0 641721
box -60594 -89821 100570 74241
use RF_switch  RF_switch_0
timestamp 1669601918
transform 0 1 535309 -1 0 212241
box -74825 -46550 34654 48242
use SCPW_M1_498p3um  SCPW_M1_498p3um_0
timestamp 1669601918
transform 0 -1 325844 1 0 294933
box -28540 -51404 28540 82036
use SCPW_M1_999p9um  SCPW_M1_999p9um_0
timestamp 1669601918
transform 0 -1 381368 1 0 142898
box -28540 -51404 28540 182356
use SCPW_M2_498um  SCPW_M2_498um_0
timestamp 1669601918
transform 0 -1 325960 1 0 372013
box -28540 -52604 28540 81976
use SCPW_M2_999um  SCPW_M2_999um_0
timestamp 1669601918
transform 0 -1 379482 1 0 215804
box -28540 -52604 28540 182176
use Standalone_mosfet_32f  Standalone_mosfet_32f_0
timestamp 1669601918
transform 0 -1 271231 1 0 56000
box -28540 -21019 32097 23598
use Standalone_mosfet_32f  Standalone_mosfet_32f_1
timestamp 1669601918
transform 0 -1 133000 1 0 216529
box -28540 -21019 32097 23598
use Standalone_mosfet_150f  Standalone_mosfet_150f_0
timestamp 1669601918
transform 0 -1 342199 1 0 56000
box -25209 -37289 31871 7178
use Standalone_mosfet_150f  Standalone_mosfet_150f_1
timestamp 1669601918
transform 0 -1 116152 1 0 139286
box -25209 -37289 31871 7178
use VGA_final  VGA_final_0
timestamp 1669601918
transform 0 1 148872 -1 0 625407
box -78593 -80722 69450 83722
use balun_v_finalstruct  balun_v_finalstruct_0
timestamp 1669601918
transform 0 -1 297697 1 0 465553
box -45000 -45000 45000 57000
use contact$2  contact$2_0
timestamp 1669601918
transform 0 -1 515842 -1 0 557834
box -320 -320 320 320
use contact$2  contact$2_1
timestamp 1669601918
transform 0 -1 509999 -1 0 557826
box -320 -320 320 320
use contact$2  contact$2_2
timestamp 1669601918
transform 1 0 10136 0 1 687958
box -320 -320 320 320
use contact$2  contact$2_3
timestamp 1669601918
transform 1 0 8330 0 1 687976
box -320 -320 320 320
use contact$2  contact$2_4
timestamp 1669601918
transform 1 0 13400 0 1 687959
box -320 -320 320 320
use contact$2  contact$2_5
timestamp 1669601918
transform 1 0 10144 0 1 684708
box -320 -320 320 320
use contact$2  contact$2_6
timestamp 1669601918
transform 1 0 13400 0 1 684708
box -320 -320 320 320
use contact$2  contact$2_7
timestamp 1669601918
transform 1 0 8330 0 1 684708
box -320 -320 320 320
use contact$4  contact$4_0
timestamp 1669601918
transform 1 0 526349 0 1 649449
box -317 -317 317 317
use contact$4  contact$4_1
timestamp 1669601918
transform 1 0 10150 0 1 682774
box -317 -317 317 317
use contact$5  contact$5_0
timestamp 1669601918
transform 1 0 44489 0 1 485342
box -423 -643 423 643
use contact$6  contact$6_0
timestamp 1669601918
transform 1 0 65216 0 1 493944
box -128 -384 128 384
use contact$6  contact$6_1
timestamp 1669601918
transform 1 0 63406 0 1 493944
box -128 -384 128 384
use contact$7  contact$7_0
timestamp 1669601918
transform 1 0 65215 0 1 493924
box -157 -397 157 397
use contact$7  contact$7_1
timestamp 1669601918
transform 1 0 63418 0 1 493924
box -157 -397 157 397
use contact$12  contact$12_0
timestamp 1669601918
transform 0 -1 575056 1 0 547972
box -7133 -6033 7133 6033
use contact$12  contact$12_1
timestamp 1669601918
transform 1 0 518026 0 1 695541
box -7133 -6033 7133 6033
use contact$14  contact$14_0
timestamp 1669601918
transform 1 0 518026 0 1 695541
box -7022 -5902 7022 5902
use contact$16  contact$16_0
timestamp 1669601918
transform 1 0 505916 0 1 415252
box -128 -64 128 64
use contact$17  contact$17_0
timestamp 1669601918
transform 1 0 505916 0 1 415252
box -157 -77 157 77
use contact$19  contact$19_0
timestamp 1669601918
transform 1 0 513831 0 1 626510
box -77 -157 77 157
use contact$19  contact$19_1
timestamp 1669601918
transform 1 0 513831 0 1 453047
box -77 -157 77 157
use contact$20  contact$20_0
timestamp 1669601918
transform 1 0 526348 0 1 597179
box -288 -288 288 288
use contact$22  contact$22_0
timestamp 1669601918
transform 1 0 515854 0 1 554615
box -384 -384 384 384
use contact$22  contact$22_1
timestamp 1669601918
transform 1 0 509967 0 1 554615
box -384 -384 384 384
use contact$22  contact$22_2
timestamp 1669601918
transform 1 0 509994 0 1 559604
box -384 -384 384 384
use contact$22  contact$22_3
timestamp 1669601918
transform 1 0 515835 0 1 559604
box -384 -384 384 384
use contact$24  contact$24_0
timestamp 1669601918
transform 1 0 509967 0 1 554615
box -533 -533 533 533
use contact$24  contact$24_1
timestamp 1669601918
transform 1 0 515854 0 1 554615
box -533 -533 533 533
use contact$24  contact$24_2
timestamp 1669601918
transform 1 0 509994 0 1 559604
box -533 -533 533 533
use contact$24  contact$24_3
timestamp 1669601918
transform 1 0 515835 0 1 559604
box -533 -533 533 533
use contact$26  contact$26_0
timestamp 1669601918
transform 1 0 515854 0 1 554615
box -437 -437 437 437
use contact$26  contact$26_1
timestamp 1669601918
transform 1 0 509967 0 1 554615
box -437 -437 437 437
use contact$26  contact$26_2
timestamp 1669601918
transform 1 0 509994 0 1 559604
box -437 -437 437 437
use contact$26  contact$26_3
timestamp 1669601918
transform 1 0 515835 0 1 559604
box -437 -437 437 437
use contact$28  contact$28_0
timestamp 1669601918
transform 1 0 509994 0 1 559604
box -622 -622 622 622
use contact$28  contact$28_1
timestamp 1669601918
transform 1 0 515835 0 1 559604
box -622 -622 622 622
use contact  contact_0
timestamp 1669601918
transform 0 -1 515812 -1 0 557864
box -397 -397 397 397
use contact  contact_1
timestamp 1669601918
transform 1 0 10106 0 1 687988
box -397 -397 397 397
use contact  contact_2
timestamp 1669601918
transform 1 0 13415 0 1 641340
box -397 -397 397 397
use contact  contact_3
timestamp 1669601918
transform 1 0 8338 0 1 557128
box -397 -397 397 397
use esd_diodes  esd_diodes_0
timestamp 1669601918
transform 0 1 10205 -1 0 690250
box 4520 -950 6580 2380
use esd_diodes  esd_diodes_1
timestamp 1669601918
transform 0 1 10205 -1 0 693497
box 4520 -950 6580 2380
use full_IC_1  full_IC_1_0
timestamp 1669601918
transform 1 0 456764 0 1 433308
box -54600 -58300 39000 93800
use out_buf  out_buf_0
timestamp 1669601918
transform 0 -1 526566 1 0 500406
box -276 -1892 10919 2293
use r_250  r_250_0
timestamp 1669602960
transform 1 0 0 0 1 0
box 513310 558091 514573 561369
use sar_adc  sar_adc_0
timestamp 1669601918
transform 0 1 45538 -1 0 493396
box 1490 0 161861 37300
use zig-zag  zig-zag_0
array 0 5 2760 0 0 0
timestamp 1669601918
transform 1 0 452127 0 1 374269
box 0 0 128 1298
use zig-zag  zig-zag_1
array 0 12 1768 0 0 0
timestamp 1669601918
transform 1 0 53502 0 1 330748
box 0 0 128 1298
<< labels >>
rlabel metal1 s 509587 556025 510407 556825 4 VDD
port 1 nsew
rlabel metal1 s 509577 556975 510407 558525 4 in
port 2 nsew
rlabel metal1 s 509567 558585 510417 558715 4 VSS
port 3 nsew
rlabel metal1 s 515433 556025 516253 556825 4 VDD
port 1 nsew
rlabel metal1 s 515423 556975 516253 558525 4 in
port 2 nsew
rlabel metal1 s 515413 558585 516263 558715 4 VSS
port 3 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 4 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 5 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 6 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 7 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 8 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 9 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 10 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 11 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 12 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 13 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 14 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 15 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 16 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 17 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 18 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 19 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 20 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 21 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 22 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 23 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 24 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 25 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 26 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 27 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 28 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 29 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 30 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 31 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 32 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 33 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 34 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 35 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 36 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 37 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 38 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 39 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 40 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 41 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 42 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 43 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 44 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 45 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 46 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 47 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 48 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 49 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 50 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 51 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 52 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 53 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 54 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 55 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 56 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 57 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 58 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 59 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 60 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 61 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 62 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 63 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 64 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 65 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 66 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 67 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 68 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 69 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 70 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 71 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 72 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 73 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 74 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 75 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 76 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 77 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 78 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 79 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 80 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 81 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 82 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 83 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 84 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 85 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 86 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 87 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 88 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 89 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 90 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 91 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 92 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 93 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 94 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 95 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 96 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 97 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 98 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 99 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 100 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 101 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 102 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 103 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 104 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 105 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 106 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 107 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 108 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 109 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 110 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 111 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 112 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 113 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 114 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 115 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 116 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 117 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 118 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 119 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 120 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 121 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 122 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 123 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 124 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 125 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 126 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 127 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 128 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 129 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 130 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 131 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 132 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 133 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 134 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 135 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 136 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 137 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 138 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 139 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 140 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 141 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 142 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 143 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 144 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 145 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 146 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 147 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 148 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 149 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 150 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 151 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 152 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 153 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 154 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 155 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 156 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 157 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 158 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 159 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 160 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 161 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 162 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 163 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 164 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 165 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 166 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 167 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 168 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 169 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 170 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 171 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 172 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 173 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 174 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 175 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 176 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 177 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 178 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 179 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 180 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 181 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 182 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 183 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 184 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 185 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 186 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 187 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 188 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 189 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 190 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 191 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 192 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 193 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 194 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 195 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 196 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 197 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 198 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 199 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 200 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 201 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 202 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 203 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 204 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 205 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 206 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 207 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 208 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 209 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 210 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 211 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 212 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 213 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 214 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 215 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 216 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 217 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 218 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 219 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 220 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 221 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 222 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 223 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 224 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 225 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 226 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 227 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 228 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 229 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 230 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 231 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 232 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 233 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 234 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 235 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 236 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 237 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 238 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 239 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 240 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 241 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 242 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 243 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 244 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 245 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 246 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 247 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 248 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 249 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 250 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 251 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 252 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 253 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 254 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 255 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 256 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 257 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 258 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 259 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 260 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 261 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 262 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 263 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 264 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 265 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 266 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 267 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 268 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 269 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 270 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 271 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 272 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 273 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 274 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 275 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 276 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 277 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 278 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 279 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 280 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 281 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 282 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 283 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 284 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 285 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 286 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 287 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 288 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 289 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 290 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 291 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 292 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 293 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 294 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 295 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 296 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 297 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 298 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 299 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 300 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 301 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 302 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 303 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 304 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 305 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 306 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 307 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 308 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 309 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 310 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 311 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 312 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 313 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 314 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 315 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 316 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 317 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 318 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 319 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 320 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 321 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 322 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 323 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 324 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 325 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 326 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 327 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 328 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 329 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 330 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 331 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 332 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 333 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 334 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 335 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 336 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 337 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 338 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 339 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 340 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 341 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 342 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 343 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 344 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 345 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 346 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 347 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 348 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 349 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 350 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 351 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 352 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 353 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 354 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 355 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 356 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 357 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 358 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 359 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 360 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 361 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 362 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 363 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 364 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 365 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 366 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 367 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 368 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 369 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 370 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 371 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 372 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 373 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 374 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 375 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 376 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 377 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 378 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 379 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 380 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 381 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 382 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 383 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 384 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 385 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 386 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 387 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 388 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 389 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 390 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 391 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 392 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 393 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 394 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 395 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 396 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 397 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 398 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 399 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 400 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 401 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 402 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 403 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 404 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 405 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 406 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 407 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 408 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 409 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 410 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 411 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 412 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 413 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 414 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 415 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 416 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 417 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 418 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 419 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 420 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 421 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 422 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 423 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 424 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 425 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 426 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 427 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 428 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 429 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 430 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 431 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 432 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 433 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 434 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 435 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 436 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 437 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 438 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 439 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 440 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 441 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 442 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 443 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 444 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 445 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 446 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 447 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 448 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 449 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 450 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 451 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 452 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 453 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 454 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 455 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 456 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 457 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 458 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 459 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 460 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 461 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 462 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 463 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 464 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 465 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 466 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 467 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 468 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 469 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 470 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 471 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 472 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 473 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 474 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 475 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 476 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 477 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 478 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 479 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 480 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 481 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 482 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 483 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 484 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 485 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 486 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 487 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 488 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 489 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 490 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 491 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 492 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 493 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 494 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 495 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 496 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 497 nsew
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 498 nsew
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 499 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 500 nsew
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 498 nsew
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 499 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 500 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 501 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 502 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 503 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 504 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 505 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 506 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 507 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 508 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 509 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 510 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 511 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 512 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 513 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 514 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 498 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 498 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 515 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 516 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 517 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 518 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 519 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 520 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 521 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 522 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 523 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 524 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 525 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 526 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 527 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 528 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 529 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 530 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 531 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 532 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 533 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 534 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 535 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 536 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 537 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 537 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 538 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 538 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 539 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 539 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 540 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 541 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 542 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 543 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 499 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 500 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 544 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 545 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 546 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 547 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 548 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 549 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 550 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 551 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 499 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 500 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 552 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 553 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 554 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 555 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 556 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 557 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 558 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 559 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 560 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 561 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 562 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 563 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 564 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 565 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 566 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 567 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 568 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 568 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 569 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 570 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 571 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 572 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 573 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 573 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 574 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 575 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 576 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 577 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 578 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 579 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 580 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 581 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 582 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 583 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 584 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 585 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 586 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 587 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 588 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 589 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 590 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 591 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 592 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 593 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 594 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 595 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 596 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 597 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 598 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 599 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 600 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 601 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 602 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 603 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 604 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 605 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 606 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 607 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 608 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 609 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 610 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 611 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 612 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 613 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 614 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 615 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 616 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 617 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 618 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 619 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 620 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 620 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 621 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 622 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 623 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 624 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 625 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 625 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 626 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 627 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 628 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 629 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 630 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 631 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 632 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 633 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 634 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 635 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 636 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 637 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 638 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 639 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 640 nsew
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 641 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 642 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 643 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 644 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 645 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 646 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 647 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 648 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 649 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 650 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 651 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 652 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 653 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 654 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 655 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 656 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 657 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 538 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 538 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 658 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 659 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 660 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 661 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 539 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 539 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 662 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 663 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 664 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 664 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 665 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 666 nsew
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 498 nsew
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 499 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 500 nsew
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 498 nsew
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 499 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 500 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string path 181.900 16033.750 1112.200 16033.750 1112.200 12112.600 1112.200 12112.600 
<< end >>
