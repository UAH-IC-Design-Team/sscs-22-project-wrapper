* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__diode_pw2nd_05v5_EUY57X a_n400_n400# a_n502_n502#
D0 a_n502_n502# a_n400_n400# sky130_fd_pr__diode_pw2nd_05v5 pj=1.6e+07u area=1.6e+13p
.ends

.subckt esd_diodes VDD in VSS dw_4600_400#
XD1 VDD in sky130_fd_pr__diode_pw2nd_05v5_EUY57X
Xsky130_fd_pr__diode_pw2nd_05v5_EUY57X_0 in VSS sky130_fd_pr__diode_pw2nd_05v5_EUY57X
.ends

.subckt VGA_final Vctrl Vgg_1v2 RF_in RF_out Vdd_1v8 Gnd
X0 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X1 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X2 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X3 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X4 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X6 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X7 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
D0 Gnd Vdd_1v8 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X8 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 Gnd RF_out sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X11 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X12 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X15 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X16 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X17 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X18 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X19 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X20 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X21 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X23 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X24 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X25 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X26 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X27 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X28 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X29 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X30 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X32 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X33 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X34 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X35 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X36 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X37 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X38 a_47_7088# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X39 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X40 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X41 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X42 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X43 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X44 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X45 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X46 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X47 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X48 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X49 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X50 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X51 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X52 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X53 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X54 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X55 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X56 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X57 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X58 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X59 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X60 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X61 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X62 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X63 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X64 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X65 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X66 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X67 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X68 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X69 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X70 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X71 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X72 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X73 Vdd_1v8 Gnd sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X74 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X75 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
R0 Vctrl a_n45858_n64215# sky130_fd_pr__res_generic_po w=2e+06u l=1.053e+07u
X76 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X77 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X78 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X79 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X80 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X81 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X82 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X83 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X84 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X85 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X86 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X87 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X88 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X89 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X90 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X91 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X92 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X93 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X94 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X95 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X96 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X97 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X98 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X99 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X100 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X101 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X102 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X103 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X104 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X105 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X106 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X107 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X108 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X109 Gnd Gnd a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X110 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X111 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X112 a_n45858_n24875# RF_in sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X113 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X114 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X115 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X116 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X117 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X118 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X119 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X120 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X121 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X122 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X123 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X124 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X125 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X126 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X127 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X128 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X129 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X130 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X131 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X132 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X133 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X134 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X135 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X136 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X137 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X138 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X139 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X140 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X141 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X142 a_n45858_n64215# Gnd sky130_fd_pr__cap_mim_m3_1 l=1.5e+07u w=1.5e+07u
X143 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X144 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X145 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X146 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X147 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X148 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X149 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X150 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X151 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X152 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X153 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X154 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X155 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X156 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X157 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X158 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X159 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X160 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X161 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X162 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X163 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X164 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X165 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X166 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X167 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X168 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X169 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X170 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X171 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X172 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X173 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X174 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X175 a_47_7088# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X176 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X177 Gnd Gnd a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X178 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X179 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X180 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X181 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X182 Gnd a_n45858_n24875# sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X183 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X184 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X185 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X186 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X187 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X188 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X189 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
D1 Gnd a_n45858_n24875# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X190 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X191 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X192 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X193 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X194 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X195 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X196 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X197 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X198 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X199 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X200 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X201 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X202 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X203 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X204 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X205 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X206 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X207 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X208 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X209 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X210 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X211 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X212 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
D2 Gnd a_n45858_n64215# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X213 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X214 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X215 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X216 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X217 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X218 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X219 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X220 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X221 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X222 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X223 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X224 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X225 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X226 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X227 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X228 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X229 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X230 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X231 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X232 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X233 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X234 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X235 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X236 Gnd RF_out sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X237 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X238 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X239 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X240 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X241 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X242 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X243 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X244 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X245 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X246 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X247 Gnd a_n45858_n24875# sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X248 Vctrl Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X249 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X250 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X251 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X252 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X253 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X254 a_n45858_n24875# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X255 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X256 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X257 a_47_7088# a_n45858_n64215# Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X258 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X259 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X260 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X261 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X262 a_n45858_n64215# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X263 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X264 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X265 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X266 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X267 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
R1 Vgg_1v2 a_n45858_n24875# sky130_fd_pr__res_generic_po w=2e+06u l=1.053e+07u
X268 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X269 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X270 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X271 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X272 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X273 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X274 a_n45858_n64215# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X275 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X276 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X277 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X278 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X279 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X280 Gnd Gnd a_n45858_n64215# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X281 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X282 Gnd Gnd Vctrl Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X283 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X284 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X285 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X286 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X287 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X288 a_47_7088# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X289 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X290 a_47_7088# a_n45858_n24875# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X291 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X292 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X293 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X294 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X295 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X296 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X297 Vdd_1v8 Vdd_1v8 a_n45858_n64215# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X298 Vdd_1v8 Vdd_1v8 Vctrl Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X299 Gnd Gnd a_n45858_n24875# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X300 Vdd_1v8 Vdd_1v8 a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X301 Vdd_1v8 a_n45858_n64215# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X302 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X303 Vctrl Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X304 Gnd a_n45858_n24875# a_47_7088# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X305 a_n45858_n24875# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X306 Vdd_1v8 Vdd_1v8 a_n45858_n24875# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_EUY57X$1 a_n400_n400# a_n502_n502#
D0 a_n502_n502# a_n400_n400# sky130_fd_pr__diode_pw2nd_05v5 pj=1.6e+07u area=1.6e+13p
.ends

.subckt esd_diodes$1 VDD in VSS dw_4600_400#
Xsky130_fd_pr__diode_pw2nd_05v5_EUY57X$1_0 in VSS sky130_fd_pr__diode_pw2nd_05v5_EUY57X$1
XD1 VDD in sky130_fd_pr__diode_pw2nd_05v5_EUY57X$1
.ends

.subckt sky130_fd_pr__res_generic_po_PL36XQ a_n200_1053# a_n200_n1483#
R0 a_n200_n1483# a_n200_1053# sky130_fd_pr__res_generic_po w=2e+06u l=1.053e+07u
.ends

.subckt r_250$1 m1_114_112# m1_112_2650# VSUBS
Xsky130_fd_pr__res_generic_po_PL36XQ_0 m1_112_2650# m1_114_112# sky130_fd_pr__res_generic_po_PL36XQ
.ends

.subckt esd vdd in dw_1628_n1498# dw_n2782_n1498# out vss
Xesd_diodes$1_0 vdd out vss dw_1628_n1498# esd_diodes$1
Xesd_diodes$1_1 vdd in vss dw_n2782_n1498# esd_diodes$1
Xr_250$1_0 out in vss r_250$1
.ends

.subckt Cascode_Amp Vgg_1v8 RF_out RF_in gnd
X0 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 gnd a_37860_8005# sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X31 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X41 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X46 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X57 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X60 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X62 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X71 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X77 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X79 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X80 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X81 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X82 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X84 gnd a_37860_8005# sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X85 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X86 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X87 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X88 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X89 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X90 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X91 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X93 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X94 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X95 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X96 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X97 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X98 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X100 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 a_38553_4766# a_37860_8005# RF_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
D0 gnd RF_in sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X102 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X103 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X104 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X105 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X106 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X107 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X108 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
D1 gnd a_37860_8005# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X109 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X110 RF_out a_37860_8005# a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X111 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X112 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X113 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 gnd RF_in a_38553_4766# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
R0 a_37860_8005# Vgg_1v8 sky130_fd_pr__res_generic_m5 w=2.532e+08u l=100000u
X117 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 a_38553_4766# RF_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X119 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X120 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X121 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_0 VPWR VGND X B A VNB VPB
X0 VPWR B a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_40_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X2 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_40_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_123_47# A a_40_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_40_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 VPWR VGND A X VNB VPB
X0 a_244_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X1 VPWR a_244_47# a_355_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=250000u
X2 X a_355_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_244_47# a_355_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
X6 X a_355_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_244_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=250000u
.ends

.subckt sky130_fd_sc_hd__dfstp_1 VPWR VGND D Q SET_B CLK VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_1 VPWR VGND B X A VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR Q RESET_B D CLK VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_1 VGND VPWR Y A VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR A X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 VGND VPWR A X VNB VPB
X0 a_283_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=500000u
X1 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_283_47# a_390_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=500000u
X3 VGND a_283_47# a_390_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X4 X a_390_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_283_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=500000u
X7 X a_390_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_1 VPWR VGND X B A VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__fa_1 VGND VPWR COUT CIN SUM A B VNB VPB
X0 a_76_199# B a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND A a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_738_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_1091_47# CIN a_995_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR CIN a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_382_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_1163_47# B a_1091_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR A a_382_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_995_47# a_76_199# a_738_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_382_413# CIN a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 SUM a_995_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_208_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VGND CIN a_738_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_76_199# B a_208_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_208_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_738_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VGND A a_1163_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_738_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_738_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_1163_413# B a_1091_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR A a_1163_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_382_47# CIN a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 a_382_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 SUM a_995_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_995_47# a_76_199# a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_76_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 a_1091_413# CIN a_995_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VGND a_76_199# COUT VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_1 VGND VPWR B Y A VNB VPB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_4 VGND VPWR Q RESET_B D CLK VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND A X VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VPWR LO HI VPB VNB
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__buf_6 VPWR VGND X A VNB VPB
X0 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_161_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A a_161_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR a_161_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_161_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_161_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VPWR A a_161_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND a_161_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 a_161_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt controller sw_n1 sw_n2 sw_n3 sw_n4 sw_n5 sw_n6 sw_n7 sw_n8 sw_n_sp1 sw_n_sp2
+ sw_n_sp3 sw_n_sp4 sw_n_sp5 sw_n_sp6 sw_n_sp7 sw_n_sp8 sw_n_sp9 sw_p1 sw_p2 sw_p3
+ sw_p4 sw_p5 sw_p6 sw_p7 sw_p8 sw_p_sp1 sw_p_sp2 sw_p_sp3 sw_p_sp4 sw_p_sp5 sw_p_sp6
+ sw_p_sp7 sw_p_sp8 sw_p_sp9 bit1 bit10 bit2 bit3 bit4 bit5 bit6 bit7 bit8 bit9 clk
+ comp_out_n comp_out_p comparator_clk done reset sw_sample VDD VSS
Xx4_x23 VDD VSS x4_x23/X x4_x23/B x4_x2/Y VSS VDD sky130_fd_sc_hd__and2_0
Xx4_x56 VDD VSS x4_x56/A x4_x56/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xx4_x78 VDD VSS x4_x79/Y x4_x78/Q fanout57/X x4_x78/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x45 VDD VSS x4_x76/A x4_x60/D x4_x6/Q VSS VDD sky130_fd_sc_hd__xor2_1
Xx4_x67 VSS VDD x4_x67/Q x4_x33/X x4_x80/D x1_x59/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x89 VSS VDD x4_x89/Y x4_x89/A VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x12 VSS VDD x4_x12/Q fanout54/X x4_x6/D x4_x95/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_26_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx1_x15 VSS VDD x1_x38/A x1_x32/D VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x37 VSS VDD x1_x37/X x1_x37/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x48 VSS VDD x1_x48/X x1_x48/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x26 VSS VDD x1_x58/A x1_x28/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x59 VSS VDD x1_x59/A x1_x59/X VSS VDD sky130_fd_sc_hd__clkbuf_2
Xx4_x84_x2 VDD VSS x4_x89/A x4_x94/X x4_x93/Q VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_5_195 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_20 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_18_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_150 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_34_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_31_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_175 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_15_32 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutput42 VDD VSS sw_p_sp1 x4_x100/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput7 VDD VSS bit2 x3_x67/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_16_197 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutput20 VDD VSS sw_n4 x4_x38/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput31 VDD VSS sw_n_sp7 x4_x69/Q VSS VDD sky130_fd_sc_hd__buf_2
Xx4_x46 VDD VSS x4_x46/X x4_x46/B x4_x1/Y VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_22_189 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx4_x35 VSS VDD x4_x35/Q x4_x26/X x4_x35/D x1_x41/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x79 VSS VDD x4_x79/Y x4_x82/A VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x57 VSS VDD x4_x57/Q fanout57/X x4_x57/D x4_x59/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x68 VSS VDD x4_x68/Q x4_x33/X x4_x68/D x1_x59/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x13 VSS VDD x4_x13/Q fanout54/X x4_x6/D x4_x98/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx1_x38 VSS VDD x1_x38/A x1_x38/X VSS VDD sky130_fd_sc_hd__clkbuf_2
Xx1_x16 VSS VDD x1_x18/A x1_x27/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x49 VSS VDD x4_x59/A x1_x49/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x27 VSS VDD x7_x27/X x1_x27/X VSS VDD sky130_fd_sc_hd__clkbuf_2
Xx4_x84_x3 VSS VDD x4_x84_x3/Y x4_x93/Q VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_8_193 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_23_32 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_23_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_177 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_18_54 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_203 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_29_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_28_184 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_162 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_176 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_44 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutput43 VDD VSS sw_p_sp2 x4_x104/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_31_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutput8 VDD VSS bit3 x3_x68/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_16_176 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_77 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput10 VDD VSS bit5 x3_x71/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput21 VDD VSS sw_n5 x4_x43/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput32 VDD VSS sw_n_sp8 x4_x71/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_30_190 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx4_x25 VSS VDD x4_x25/Q x4_x23/X x4_x4/D x1_x38/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_22_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x58 VSS VDD x4_x59/X x4_x58/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xx4_x69 VSS VDD x4_x69/Q x4_x36/X x4_x80/D x1_x59/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x36 VDD VSS x4_x36/X x4_x36/B x4_x89/Y VSS VDD sky130_fd_sc_hd__and2_0
Xx4_x14 VSS VDD x4_x14/Q fanout54/X x4_x6/D x1_x69/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x47 VDD VSS x4_x47/X x4_x47/B x4_x90/Y VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_26_43 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx3_x80 VSS VDD x3_x80/Q fanout71/X x3_x80/D x3_x82/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_13_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx1_x39 VSS VDD x4_x50/A x1_x62/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x17 VSS VDD x1_x17/X x1_x18/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x28 VSS VDD x7_x27/X x1_x28/X VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_8_161 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx2 VDD VSS x2/X x2/B x6/Y VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_2_189 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_22_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_119 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput44 VDD VSS sw_p_sp3 x4_x35/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_31_33 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutput9 VDD VSS bit4 x3_x70/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_16_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput11 VDD VSS bit6 x3_x74/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput22 VDD VSS sw_n6 x4_x75/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput33 VDD VSS sw_n_sp9 x4_x61/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_31_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x48 VSS VDD x4_x48/Q x4_x46/B x4_x48/D x4_x50/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x37 VDD VSS x4_x82/A x4_x54/D x4_x6/Q VSS VDD sky130_fd_sc_hd__xor2_1
Xx4_x26 VDD VSS x4_x26/X x4_x46/B x4_x26/A VSS VDD sky130_fd_sc_hd__and2_0
Xx4_x59 VDD VSS x4_x59/A x4_x59/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xx4_x15 VSS VDD x4_x15/Q fanout54/X x4_x6/D x1_x75/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_26_55 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx3_x70 VSS VDD x3_x70/Q x2/B x3_x70/D x1_x76/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_13_169 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_13_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_7_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx3_x81 VSS VDD x3_x81/Q x2/B x4_x15/Q x3_x82/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_9_118 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx1_x18 VSS VDD x1_x18/X x1_x18/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x29 VSS VDD x1_x29/X x1_x29/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_8_173 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_124 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_29_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_28_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_68 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_6_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_120 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xoutput34 VDD VSS sw_p1 x4_x22/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput45 VDD VSS sw_p_sp4 x4_x108/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_31_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_25_123 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_15_57 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutput23 VDD VSS sw_n7 x4_x77/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput12 VDD VSS bit7 x3_x75/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_31_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x49 VSS VDD x4_x50/X x4_x49/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xx4_x27 VSS VDD x4_x27/Q x4_x26/X x4_x8/D x1_x41/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x16 VDD VSS x4_x16/X x4_x46/B x4_x19/Y VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_11_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x38 VDD VSS x4_x76/A x4_x38/Q fanout54/X x4_x38/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx3_x82 VSS VDD x3_x82/Y x3_x82/A VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_26_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx3_x71 VSS VDD x3_x71/Q x2/B x3_x71/D x3_x82/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx1_x19 VSS VDD x1_x19/X x1_x29/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_21_181 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_13_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_185 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_100 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput35 VDD VSS sw_p2 x4_x106/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput46 VDD VSS sw_p_sp5 x4_x112/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_31_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_25_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx7_x14 VSS VDD x7_x19/A x7_x9/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xoutput24 VDD VSS sw_n8 x4_x80/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput13 VDD VSS bit8 x3_x78/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_31_149 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_22_116 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x17 VDD VSS x4_x17/X x4_x17/B x4_x20/Y VSS VDD sky130_fd_sc_hd__and2_0
Xx4_x28 VDD VSS x4_x6/D x4_x28/Q fanout54/X x4_x28/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx3_x72 VSS VDD x3_x69/CIN x3_x72/CIN x3_x74/D x4_x9/Q x4_x6/Q VSS VDD sky130_fd_sc_hd__fa_1
XFILLER_13_149 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_3_28 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_153 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_12_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xfanout70 VSS VDD x2/B fanout72/X VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx1_x1 VSS VDD x1_x2/D fanout60/X x1_x1/D x1_x19/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x30_x1 VDD VSS x4_x28/CLK x4_x52/X x4_x30_x3/Y VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_1_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_47 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_79 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_25_147 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx7_x26 VSS VDD x7_x27/A x7_x26/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xoutput36 VDD VSS sw_p3 x4_x114/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput47 VDD VSS sw_p_sp6 x4_x68/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_16_114 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutput25 VDD VSS sw_n_sp1 x4_x102/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput14 VDD VSS bit9 x3_x79/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_30_183 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x29 VDD VSS x4_x8/D x4_x48/D x4_x3/Q VSS VDD sky130_fd_sc_hd__xor2_1
Xx4_x18 VSS VDD x4_x26/A x4_x18/A VSS VDD sky130_fd_sc_hd__inv_1
XPHY_0 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_36 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx3_x62 VSS VDD x3_x80/D x3_x62/CIN x3_x67/D x4_x4/Q x4_x3/Q VSS VDD sky130_fd_sc_hd__fa_1
XFILLER_13_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx3_x73 VSS VDD x3_x72/CIN x3_x73/CIN x3_x75/D x4_x11/Q x4_x64/A VSS VDD sky130_fd_sc_hd__fa_1
XFILLER_12_172 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x1 VSS VDD x4_x1/Y x4_x1/A VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_12_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx6 VSS VDD x6/B x6/Y x6/A VSS VDD sky130_fd_sc_hd__xnor2_1
XFILLER_5_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_190 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xfanout71 VSS VDD fanout72/X fanout71/X VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout60 VSS VDD fanout60/X fanout61/X VSS VDD sky130_fd_sc_hd__clkbuf_4
Xx4_x30_x2 VDD VSS x4_x2/A x4_x52/X x4_x51/Q VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_34_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx1_x2 VSS VDD x1_x3/D fanout60/X x1_x2/D x1_x29/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_19_156 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_25_159 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx7_x27 VSS VDD x7_x27/X x7_x27/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xoutput37 VDD VSS sw_p4 x4_x116/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput48 VDD VSS sw_p_sp7 x4_x70/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_33_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_192 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_126 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx7_x1 VDD VSS x7_x1/A x7_x4/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput15 VDD VSS comparator_clk x5_x25/X VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_0_203 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xoutput26 VDD VSS sw_n_sp2 x4_x25/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_30_162 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x19 VSS VDD x4_x19/Y x4_x19/A VSS VDD sky130_fd_sc_hd__inv_1
XPHY_1 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx3_x74 VSS VDD x3_x74/Q x2/B x3_x74/D x3_x82/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x2 VSS VDD x4_x2/Y x4_x2/A VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_5_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx4_x44_x1 VDD VSS x4_x43/CLK x4_x63/X x4_x44_x3/Y VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_23_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xfanout72 VSS VDD input4/X fanout72/X VSS VDD sky130_fd_sc_hd__clkbuf_2
Xx4_x30_x3 VSS VDD x4_x30_x3/Y x4_x51/Q VSS VDD sky130_fd_sc_hd__inv_1
Xfanout61 VDD VSS fanout61/X x1_x37/X VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_1_161 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_34_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx1_x3 VSS VDD x1_x4/D fanout60/X x1_x3/D x1_x30/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x39_x1 VDD VSS x4_x38/CLK x4_x58/X x4_x39_x3/Y VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_3_201 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx7_x17 VDD VSS x7_x3/X x7_x1/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput38 VDD VSS sw_p5 x4_x118/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput49 VDD VSS sw_p_sp8 x4_x72/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput16 VDD VSS done x3_x82/Y VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_33_160 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx7_x2 VDD VSS x7_x2/B x7_x3/A x26/A VSS VDD sky130_fd_sc_hd__xor2_1
Xoutput27 VDD VSS sw_n_sp3 x4_x27/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_31_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_2 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_26_16 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx3_x64 VSS VDD x3_x62/CIN x3_x64/CIN x3_x68/D x4_x5/Q x4_x3/Q VSS VDD sky130_fd_sc_hd__fa_1
Xx3_x75 VSS VDD x3_x75/Q x2/B x3_x75/D x3_x82/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_32_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_12_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x3 VSS VDD x4_x3/Q x4_x23/B x4_x4/D x1_x38/X VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_12_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_159 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_17_200 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x44_x2 VDD VSS x4_x20/A x4_x63/X x4_x60/Q VSS VDD sky130_fd_sc_hd__and2_0
Xfanout73 VSS VDD input1/X x5_x28/A VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout62 VDD VSS x4_x80/D x4_x76/A VSS VDD sky130_fd_sc_hd__buf_2
Xx4_x39_x2 VDD VSS x4_x19/A x4_x58/X x4_x57/Q VSS VDD sky130_fd_sc_hd__and2_0
Xx1_x4 VSS VDD x1_x5/D fanout60/X x1_x4/D x1_x33/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_20_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_1_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_29_16 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_32_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xoutput39 VDD VSS sw_p6 x4_x74/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_25_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx7_x3 VDD VSS x7_x3/A x7_x3/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput17 VDD VSS sw_n1 x4_x21/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput28 VDD VSS sw_n_sp4 x4_x41/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_24_172 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_106 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx3_x65 VSS VDD x3_x64/CIN x3_x65/CIN x3_x70/D x4_x7/Q x4_x6/Q VSS VDD sky130_fd_sc_hd__fa_1
XPHY_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_74 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx3_x76 VSS VDD x3_x73/CIN x3_x76/CIN x3_x78/D x4_x12/Q x4_x64/A VSS VDD sky130_fd_sc_hd__fa_1
XFILLER_12_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x4 VSS VDD x4_x4/Q x4_x23/B x4_x4/D x4_x50/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_32_204 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx4_x44_x3 VSS VDD x4_x44_x3/Y x4_x60/Q VSS VDD sky130_fd_sc_hd__inv_1
Xfanout74 VDD VSS input1/X x5_x19/CLK VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout63 VDD VSS x4_x76/A x4_x9/D VSS VDD sky130_fd_sc_hd__buf_2
Xfanout52 VSS VDD x4_x36/B x4_x47/B VSS VDD sky130_fd_sc_hd__clkbuf_4
Xx1_x5 VSS VDD x1_x6/D fanout61/X x1_x5/D x1_x47/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_18_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x39_x3 VSS VDD x4_x39_x3/Y x4_x57/Q VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_24_72 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_29_28 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_96 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx7_x19 VSS VDD x7_x26/A x7_x19/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx7_x4 VDD VSS x7_x4/A x7_x5/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xoutput18 VDD VSS sw_n2 x4_x28/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput29 VDD VSS sw_n_sp5 x4_x110/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_21_84 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_21_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_15_184 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_4 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx3_x77 VSS VDD x3_x76/CIN x4_x14/Q x3_x79/D x4_x13/Q x4_x64/A VSS VDD sky130_fd_sc_hd__fa_1
XFILLER_8_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x5 VSS VDD x4_x5/Q x4_x46/B x4_x8/D x4_x53/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_7_191 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_27_94 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_43 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xfanout64 VDD VSS x4_x6/D x4_x9/D VSS VDD sky130_fd_sc_hd__buf_2
Xfanout53 VSS VDD x4_x17/B x4_x47/B VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_13_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx1_x6 VSS VDD x1_x7/D fanout60/X x1_x6/D x1_x48/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_34_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_138 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_18_193 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx7_x5 VDD VSS x7_x5/A x7_x6/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_24_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xoutput19 VDD VSS sw_n3 x4_x32/Q VSS VDD sky130_fd_sc_hd__buf_2
XPHY_5 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx3_x67 VSS VDD x3_x67/Q x2/B x3_x67/D x3_x82/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_21_144 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx3_x78 VSS VDD x3_x78/Q x2/B x3_x78/D x3_x82/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_35_203 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_32_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_16_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx4_x6 VSS VDD x4_x6/Q fanout54/X x4_x6/D x1_x41/X VSS VDD sky130_fd_sc_hd__dfrtp_4
XFILLER_4_77 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_4_99 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xfanout65 VDD VSS x4_x4/D x4_x8/D VSS VDD sky130_fd_sc_hd__buf_2
Xfanout54 VSS VDD fanout54/X x4_x17/B VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_13_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx4_x85_x1 VDD VSS x4_x81/CLK x4_x97/X x4_x85_x3/Y VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_1_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx1_x7 VSS VDD x1_x8/D fanout60/X x1_x7/D x1_x51/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_34_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_24_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx7_x6 VDD VSS x7_x6/A x7_x9/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_24_197 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_6 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_30_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx3_x68 VSS VDD x3_x68/Q x2/B x3_x68/D x3_x82/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_21_156 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx3_x79 VSS VDD x3_x79/Q x2/B x3_x79/D x3_x82/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_7_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_32_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_32_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_16_97 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_75 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_189 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx4_x7 VSS VDD x4_x7/Q x4_x46/B x4_x8/D x4_x56/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_4_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xfanout55 VSS VDD x4_x46/B fanout57/X VSS VDD sky130_fd_sc_hd__clkbuf_4
Xx4_x85_x2 VDD VSS x4_x90/A x4_x97/X x4_x96/Q VSS VDD sky130_fd_sc_hd__and2_0
Xfanout66 VDD VSS x4_x8/D x4_x82/A VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_13_65 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx1_x8 VSS VDD x1_x9/D fanout60/X x1_x8/D x1_x52/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_24_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_1_79 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xinput1 VSS VDD input1/X clk VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_19_31 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_35_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_19_86 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_173 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_7 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx3_x69 VSS VDD x3_x65/CIN x3_x69/CIN x3_x71/D x4_x8/Q x4_x6/Q VSS VDD sky130_fd_sc_hd__fa_1
XFILLER_32_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_29_202 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_179 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x8 VSS VDD x4_x8/Q x4_x46/B x4_x8/D x4_x59/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_27_75 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_197 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x85_x3 VSS VDD x4_x85_x3/Y x4_x96/Q VSS VDD sky130_fd_sc_hd__inv_1
Xfanout56 VSS VDD fanout57/X x4_x23/B VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout67 VDD VSS x4_x82/A x4_x9/D VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_13_77 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx1_x9 VSS VDD x1_x9/Q fanout60/X x1_x9/D x1_x53/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_24_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_65 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xinput2 VSS VDD x7_x2/B comp_out_n VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_35_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_174 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_21_33 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_30_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_8 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_21_169 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_11_191 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x9 VSS VDD x4_x9/Q x4_x17/B x4_x9/D x4_x86/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_27_87 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_32 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xfanout68 VSS VDD x25/X x4_x9/D VSS VDD sky130_fd_sc_hd__clkbuf_2
Xfanout57 VSS VDD fanout57/X x4_x17/B VSS VDD sky130_fd_sc_hd__clkbuf_4
XFILLER_1_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_24_11 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xinput3 VSS VDD x26/A comp_out_p VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_27_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx7_x9 VSS VDD x7_x9/X x7_x9/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_24_123 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_30_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_15_101 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_21_104 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_44 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_90 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_4_111 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_166 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xfanout69 VSS VDD x1_x35/B fanout72/X VSS VDD sky130_fd_sc_hd__clkbuf_4
Xfanout58 VDD VSS x28/X x4_x17/B VSS VDD sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_57 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_13_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_1_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_5_91 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_23 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_202 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_6_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xinput4 VSS VDD input4/X reset VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_27_121 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_19_12 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_47 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_10_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_18_8 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_24_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_15_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_15 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_7_142 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_4_123 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_4_178 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xfanout59 VSS VDD x1_x76/X x3_x82/A VSS VDD sky130_fd_sc_hd__clkbuf_2
XFILLER_1_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_1_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_19_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_136 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_21_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_15_169 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_7_38 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_68 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_81 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_4_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_1_149 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_35_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_35_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_170 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_181 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_15_159 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_23_8 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_21_118 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_16_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_151 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_27_25 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_4_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x34_x1 VDD VSS x4_x32/CLK x4_x55/X x4_x34_x3/Y VSS VDD sky130_fd_sc_hd__and2_0
Xx5_x1 VSS VDD x5_x1/X x5_x1/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_0_183 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_14_92 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_18_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_24_149 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_16_8 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_108 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx5_x2 VSS VDD x5_x3/A x5_x4/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx4_x34_x2 VDD VSS x4_x18/A x4_x55/X x4_x54/Q VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_19_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_10_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_70 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_18_147 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_2_63 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_11_72 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_16_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_20_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_120 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx1_x36_75 VSS VDD x1_x36_75/LO x1_x36/A VDD VSS sky130_fd_sc_hd__conb_1
Xx5_x3 VDD VSS x5_x3/X x5_x3/A VSS VDD sky130_fd_sc_hd__buf_6
Xx4_x34_x3 VSS VDD x4_x34_x3/Y x4_x54/Q VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_12_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_5_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_71 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_33_107 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_60 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_2_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_20_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x132 VSS VDD x4_x132/Q fanout57/X x4_x133/Y x1_x69/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_21_8 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x110 VSS VDD x4_x110/Q x4_x17/X x4_x9/D x1_x41/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_11_198 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx5_x4 VSS VDD x5_x4/X x5_x7/D VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_3_161 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_71 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_24_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_14_73 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_27_127 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_50 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_32_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx5_x20 VSS VDD x5_x21/D x1_x35/B x5_x20/D x5_x28/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_14_163 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_11_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_11_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_35_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_32_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x100 VSS VDD x4_x100/Q x4_x46/X x4_x99/Y x1_x38/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x133 VSS VDD x4_x133/Y x4_x82/A VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x111 VSS VDD x4_x111/Y x4_x8/D VSS VDD sky130_fd_sc_hd__inv_1
Xx30 VSS VDD x30/X x30/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_11_144 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_31_206 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx5_x5 VSS VDD x5_x7/D x1_x35/B x5_x5/D x5_x28/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_28_94 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_30_51 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_85 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_41 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_27_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_19 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_35_183 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_35_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_27_139 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_62 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_51 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx5_x21 VSS VDD x5_x22/A x1_x35/B x5_x21/D x5_x28/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx5_x10 VSS VDD x5_x11/D x1_x35/B x5_x9/Q x5_x28/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_15_109 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx4_x83_x1 VDD VSS x4_x75/CLK x4_x91/X x4_x83_x3/Y VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_14_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_14_175 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_11_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_32_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_28_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx4_x112 VSS VDD x4_x112/Q x4_x17/X x4_x113/Y x1_x41/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_8_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_8_98 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_33_95 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_63 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx5_x6 VDD VSS x5_x6/A x5_x6/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_155 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_10_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_53 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_30_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_35_162 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_63 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_52 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_74 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_18_107 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XPHY_30 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx5_x22 VSS VDD x5_x5/D x5_x22/A VSS VDD sky130_fd_sc_hd__inv_1
Xx5_x11 VSS VDD x5_x12/D x1_x35/B x5_x11/D x5_x28/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x83_x2 VDD VSS x4_x88/A x4_x91/X x4_x87/Q VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_23_121 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_23_143 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_135 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x102 VSS VDD x4_x102/Q x4_x46/X x4_x4/D x1_x38/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_22_75 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_22_42 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x113 VSS VDD x4_x113/Y x4_x8/D VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_11_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_7_106 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_75 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx5_x7 VSS VDD x5_x8/D x1_x35/B x5_x7/D x5_x28/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_28_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_28_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_45 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_14_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_30_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_64 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_53 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_42 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_31 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx4_x83_x3 VSS VDD x4_x83_x3/Y x4_x87/Q VSS VDD sky130_fd_sc_hd__inv_1
Xx5_x12 VSS VDD x5_x13/D x1_x35/B x5_x12/D x5_x28/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx5_x23 VDD VSS x5_x1/A x5_x24/Y x5_x6/X VSS VDD sky130_fd_sc_hd__and2_1
XFILLER_23_155 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_23_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_14_122 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x103 VSS VDD x4_x104/D x4_x4/D VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x114 VDD VSS x4_x115/Y x4_x114/Q x4_x46/B x4_x32/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx1_x70 VSS VDD x1_x70/X x1_x3/D VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_11_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_11_158 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_8_34 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_98 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_87 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx5_x8 VSS VDD x5_x9/D x1_x35/B x5_x8/D x5_x28/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_35_175 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_65 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_54 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_32 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_21 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_10 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx5_x13 VSS VDD x5_x14/D fanout72/X x5_x13/D x5_x19/CLK VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx5_x24 VSS VDD x5_x24/Y x5_x3/X VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_14_134 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx4_x90 VSS VDD x4_x90/Y x4_x90/A VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x104 VSS VDD x4_x104/Q x4_x23/X x4_x104/D x1_x38/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x115 VSS VDD x4_x115/Y x4_x4/D VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_22_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx1_x60 VSS VDD x1_x65/A x1_x8/D VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x71 VSS VDD x1_x75/A x1_x71/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_26_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_10_170 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_33_43 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx5_x9 VSS VDD x5_x9/Q x1_x35/B x5_x9/D x5_x28/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_0_147 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_0_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_66 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_55 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_187 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_25_99 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_44 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_33 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_22 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_11 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx5_x14 VSS VDD x5_x15/D fanout72/X x5_x14/D x5_x19/CLK VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_23_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx5_x25 VSS VDD x5_x25/X x5_x27/X VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_14_113 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x80 VDD VSS x4_x80/D x4_x80/Q x4_x36/B x4_x81/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x91 VSS VDD x4_x92/X x4_x91/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xx4_x105 VSS VDD x4_x22/D x4_x4/D VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x116 VDD VSS x4_x117/Y x4_x116/Q x4_x46/B x4_x38/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx1_x50 VSS VDD x4_x86/A x1_x50/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x72 VSS VDD x1_x76/A x1_x72/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x61 VSS VDD x1_x67/A x1_x9/D VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_19_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_6_197 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_8_69 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_0_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_5_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_14_79 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_155 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_12 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_67 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_56 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_67 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_45 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_188 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_34 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_23 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx5_x15 VSS VDD x5_x16/D fanout72/X x5_x15/D x5_x19/CLK VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_23_169 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_23_103 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx5_x26 VSS VDD x5_x27/A x5_x1/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx4_x81 VDD VSS x4_x82/Y x4_x81/Q fanout57/X x4_x81/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x70 VSS VDD x4_x70/Q x4_x36/X x4_x70/D x1_x59/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_2_9 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x92 VDD VSS x4_x92/A x4_x92/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_20_128 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_9_184 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x106 VDD VSS x4_x107/Y x4_x106/Q x4_x23/B x4_x28/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x117 VSS VDD x4_x117/Y x4_x82/A VSS VDD sky130_fd_sc_hd__inv_1
Xx1_x62 VSS VDD x1_x62/X x1_x1/D VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x40 VSS VDD x4_x53/A x1_x66/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx25 VSS VDD x25/X x27/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x73 VSS VDD x1_x77/A x1_x73/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x51 VSS VDD x1_x51/X x1_x52/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_6_121 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_3_113 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_31_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_5_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_14_14 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_68 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_46 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_35 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_24 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_39 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_2_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_1_200 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_13 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx5_x16 VSS VDD x5_x17/D fanout71/X x5_x16/D x5_x19/CLK VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx5_x27 VSS VDD x5_x27/X x5_x27/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_31_181 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x82 VSS VDD x4_x82/Y x4_x82/A VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x60 VSS VDD x4_x60/Q x4_x47/B x4_x60/D x4_x86/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_14_104 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x71 VSS VDD x4_x71/Q x4_x47/X x4_x80/D x1_x59/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x93 VSS VDD x4_x93/Q x4_x36/B x4_x93/D x4_x95/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_9_130 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_9_152 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x107 VSS VDD x4_x107/Y x4_x4/D VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x118 VDD VSS x4_x119/Y x4_x118/Q fanout57/X x4_x43/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx1_x41 VSS VDD x1_x70/X x1_x41/X VSS VDD sky130_fd_sc_hd__clkbuf_2
Xx1_x30 VSS VDD x1_x30/X x1_x33/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx26 VSS VDD x27/A x26/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x52 VSS VDD x1_x52/X x1_x52/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x63 VSS VDD x1_x68/A x1_x9/Q VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x74 VSS VDD x1_x78/A x1_x74/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_6_133 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_33_57 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_3_169 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_24_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x24_x1 VDD VSS x4_x22/CLK x4_x49/X x4_x24_x3/Y VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_28_24 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_176 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_29_165 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_35_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_20_80 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_60 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_69 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_34_190 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_58 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_26_124 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_47 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_36 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_25 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_14 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_32_105 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_113 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xx5_x17 VSS VDD x5_x18/D fanout71/X x5_x17/D x5_x19/CLK VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx5_x28 VDD VSS x5_x28/A x5_x6/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xx4_x50 VDD VSS x4_x50/A x4_x50/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xx4_x72 VSS VDD x4_x72/Q x4_x47/X x4_x73/Y x1_x59/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x61 VSS VDD x4_x61/Q x4_x36/B x4_x80/D x1_x69/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x94 VSS VDD x4_x95/X x4_x94/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xx4_x119 VSS VDD x4_x119/Y x4_x82/A VSS VDD sky130_fd_sc_hd__inv_1
Xx1_x31 VSS VDD x1_x32/D fanout60/X x1_x36/X x1_x17/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx1_x20 VSS VDD x1_x29/A x1_x27/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx4_x108 VSS VDD x4_x108/Q x4_x16/X x4_x111/Y x1_x41/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx1_x42 VSS VDD x1_x46/A x1_x4/D VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx27 VSS VDD x27/X x27/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x53 VSS VDD x1_x53/X x1_x54/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x64 VSS VDD x1_x69/A x1_x64/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x75 VSS VDD x1_x75/X x1_x75/A VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_9_142 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_9_164 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_33_200 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_12_70 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_163 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_167 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_17_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_3_137 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x24_x2 VDD VSS x4_x1/A x4_x49/X x4_x48/Q VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_17_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_203 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_30_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_30_15 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_35_147 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_125 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_59 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_26 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_48 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_37 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_26 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_15 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_32_128 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_17_169 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx5_x18 VSS VDD x5_x19/D fanout71/X x5_x18/D x5_x19/CLK VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_31_161 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_11_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xx4_x51 VSS VDD x4_x51/Q x4_x46/B x4_x51/D x4_x53/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x40 VDD VSS x4_x82/A x4_x57/D x4_x6/Q VSS VDD sky130_fd_sc_hd__xor2_1
Xx4_x62 VDD VSS x4_x80/D x4_x93/D x4_x64/A VSS VDD sky130_fd_sc_hd__xor2_1
Xx4_x95 VDD VSS x4_x95/A x4_x95/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xx4_x73 VSS VDD x4_x73/Y x4_x76/A VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_20_109 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx28 VSS VDD x28/X x30/X VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_13_161 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_40 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_3_62 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx1_x32 VSS VDD x1_x1/D fanout60/X x1_x32/D x1_x18/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x109 VSS VDD x4_x35/D x4_x8/D VSS VDD sky130_fd_sc_hd__inv_1
Xx1_x21 VSS VDD x1_x33/A x1_x27/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x43 VSS VDD x1_x49/A x1_x5/D VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x54 VSS VDD x1_x54/X x1_x54/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x76 VSS VDD x1_x76/X x1_x76/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x65 VSS VDD x4_x92/A x1_x65/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x10 VSS VDD x1_x64/A fanout61/X x1_x9/Q x1_x54/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_33_9 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_10_131 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_149 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x24_x3 VSS VDD x4_x24_x3/Y x4_x48/Q VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_0_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_0_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_35_137 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_25_38 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_49 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_38 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_27 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_6_51 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_6_95 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_16 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_17_159 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx5_x19 VSS VDD x5_x20/D fanout71/X x5_x19/D x5_x19/CLK VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x52 VSS VDD x4_x53/X x4_x52/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xx4_x41 VSS VDD x4_x41/Q x4_x16/X x4_x6/D x1_x41/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x63 VSS VDD x4_x86/X x4_x63/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xx4_x74 VDD VSS x4_x76/Y x4_x74/Q x4_x47/B x4_x75/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
XFILLER_7_3 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x96 VSS VDD x4_x96/Q x4_x36/B x4_x96/D x4_x98/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx29 VSS VDD x30/A x2/X VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_13_184 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_3_52 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx1_x66 VSS VDD x1_x66/X x1_x2/D VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x33 VSS VDD x1_x33/X x1_x33/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x22 VSS VDD x1_x48/A x1_x27/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x44 VSS VDD x1_x50/A x1_x6/D VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x55 VSS VDD x1_x55/X x1_x56/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x77 VSS VDD x6/A x1_x77/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x11 VSS VDD x1_x71/A fanout61/X x1_x64/A x1_x55/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_3_96 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_0_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_40 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_9_84 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_18_71 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_22_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_14_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XPHY_28 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_17 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_39 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_31_174 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xx4_x31 VDD VSS x4_x4/D x4_x51/D x4_x3/Q VSS VDD sky130_fd_sc_hd__xor2_1
Xx4_x53 VDD VSS x4_x53/A x4_x53/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_22_163 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x20 VSS VDD x4_x20/Y x4_x20/A VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x86 VDD VSS x4_x86/A x4_x86/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
Xx4_x75 VDD VSS x4_x80/D x4_x75/Q x4_x36/B x4_x75/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x64 VDD VSS x4_x80/D x4_x96/D x4_x64/A VSS VDD sky130_fd_sc_hd__xor2_1
Xx4_x42 VDD VSS x4_x76/A x4_x87/D x4_x64/A VSS VDD sky130_fd_sc_hd__xor2_1
Xx4_x97 VSS VDD x4_x98/X x4_x97/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xx1_x34 VSS VDD x1_x35/A x5_x3/X VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_22_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx1_x45 VSS VDD x1_x59/A x1_x7/D VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x23 VSS VDD x1_x52/A x1_x28/X VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x78 VSS VDD x6/B x1_x78/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x56 VSS VDD x1_x56/X x1_x56/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x67 VSS VDD x4_x95/A x1_x67/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x12 VSS VDD x1_x72/A fanout61/X x1_x71/A x1_x56/X VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_10_177 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_17_29 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_28_17 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_34_60 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_18_61 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_34_183 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_26_117 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XPHY_29 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XPHY_18 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xoutput50 VDD VSS sw_p_sp9 x4_x132/Q VSS VDD sky130_fd_sc_hd__buf_2
Xx4_x54 VSS VDD x4_x54/Q fanout57/X x4_x54/D x4_x56/A VSS VDD sky130_fd_sc_hd__dfrtp_1
XFILLER_16_183 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx4_x76 VSS VDD x4_x76/Y x4_x76/A VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x21 VDD VSS x4_x6/D x4_x21/Q fanout54/X x4_x22/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x32 VDD VSS x4_x6/D x4_x32/Q fanout54/X x4_x32/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x65 VSS VDD x4_x68/D x4_x76/A VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x43 VDD VSS x4_x76/A x4_x43/Q x4_x36/B x4_x43/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x87 VSS VDD x4_x87/Q x4_x36/B x4_x87/D x4_x92/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x10 VSS VDD x4_x64/A x4_x47/B x4_x80/D x1_x59/X VSS VDD sky130_fd_sc_hd__dfrtp_4
Xx4_x98 VDD VSS x4_x98/A x4_x98/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_22_197 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
Xx1_x35 VDD VSS x1_x37/A x1_x35/B x1_x35/A VSS VDD sky130_fd_sc_hd__and2_1
Xx1_x46 VSS VDD x4_x56/A x1_x46/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x13 VSS VDD x1_x73/A fanout61/X x1_x72/A x1_x57/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx1_x57 VSS VDD x1_x57/X x1_x58/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x68 VSS VDD x4_x98/A x1_x68/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x24 VSS VDD x1_x54/A x1_x28/X VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_12_96 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_12_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_12_63 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_10_189 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_3_108 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_73 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_2_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_28_29 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_18_40 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_29_126 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_85 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_41 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_19_181 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XPHY_19 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
Xoutput40 VDD VSS sw_p7 x4_x78/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput51 VDD VSS sw_sample x5_x3/X VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_31_84 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput5 VDD VSS bit1 x3_x80/Q VSS VDD sky130_fd_sc_hd__buf_2
Xx4_x22 VDD VSS x4_x22/D x4_x22/Q x4_x23/B x4_x22/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x33 VDD VSS x4_x33/X x4_x36/B x4_x88/Y VSS VDD sky130_fd_sc_hd__and2_0
Xx4_x11 VSS VDD x4_x11/Q fanout54/X x4_x6/D x4_x92/A VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx4_x99 VSS VDD x4_x99/Y x4_x4/D VSS VDD sky130_fd_sc_hd__inv_1
XFILLER_22_132 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x55 VSS VDD x4_x56/X x4_x55/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xx4_x77 VDD VSS x4_x80/D x4_x77/Q x4_x36/B x4_x78/CLK VSS VDD sky130_fd_sc_hd__dfstp_1
Xx4_x88 VSS VDD x4_x88/Y x4_x88/A VSS VDD sky130_fd_sc_hd__inv_1
Xx4_x66 VSS VDD x4_x70/D x4_x76/A VSS VDD sky130_fd_sc_hd__inv_1
Xx1_x36 VSS VDD x1_x36/X x1_x36/A VSS VDD sky130_fd_sc_hd__buf_1
Xx1_x47 VSS VDD x1_x47/X x1_x48/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x69 VDD VSS x1_x69/X x1_x69/A VSS VDD sky130_fd_sc_hd__buf_2
Xx1_x14 VSS VDD x1_x74/A fanout61/X x1_x73/A x1_x58/X VSS VDD sky130_fd_sc_hd__dfrtp_1
Xx1_x58 VSS VDD x1_x58/X x1_x58/A VSS VDD sky130_fd_sc_hd__clkbuf_1
Xx1_x25 VSS VDD x1_x56/A x1_x28/X VSS VDD sky130_fd_sc_hd__clkbuf_1
XFILLER_9_169 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_27_202 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
Xx4_x84_x1 VDD VSS x4_x78/CLK x4_x94/X x4_x84_x3/Y VSS VDD sky130_fd_sc_hd__and2_0
XFILLER_10_124 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_5_3 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_33_19 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_96 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
XFILLER_23_85 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_153 VDD VSS VSS VDD sky130_fd_sc_hd__decap_3
XFILLER_2_197 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_29_138 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_20_97 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
XFILLER_20_20 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_34_141 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_20_3 VDD VSS VSS VDD sky130_fd_sc_hd__decap_6
Xoutput41 VDD VSS sw_p8 x4_x81/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_25_130 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
XFILLER_17_119 VSS VDD VSS VDD sky130_ef_sc_hd__decap_12
XFILLER_15_20 VSS VDD VSS VDD sky130_fd_sc_hd__decap_4
Xoutput6 VDD VSS bit10 x3_x81/Q VSS VDD sky130_fd_sc_hd__buf_2
Xoutput30 VDD VSS sw_n_sp6 x4_x67/Q VSS VDD sky130_fd_sc_hd__buf_2
XFILLER_16_141 VDD VSS VSS VDD sky130_fd_sc_hd__decap_8
.ends

.subckt sky130_fd_pr__nfet_01v8_9CGS2F a_n33_n148# a_15_n60# a_n73_n60# VSUBS
X0 a_15_n60# a_n33_n148# a_n73_n60# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_46WN3R a_n73_n129# a_n33_n226# a_15_n129# w_n109_n229#
X0 a_15_n129# a_n33_n226# a_n73_n129# w_n109_n229# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_5XXJZ8 a_n33_n91# a_n105_n179# a_63_n91# a_n125_n91#
+ VSUBS
X0 a_63_n91# a_n105_n179# a_n33_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X1 a_n33_n91# a_n105_n179# a_n125_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_CBMBZG a_n33_n165# a_n125_n165# w_n169_n265# a_63_n165#
+ a_n85_n262#
X0 a_n33_n165# a_n85_n262# a_n125_n165# w_n169_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X1 a_63_n165# a_n85_n262# a_n33_n165# w_n169_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ZDVJZL a_159_n91# a_n221_n91# a_n33_n91# a_n179_n179#
+ a_63_n91# a_n129_n91# VSUBS
X0 a_63_n91# a_n179_n179# a_n33_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X1 a_n33_n91# a_n179_n179# a_n129_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X2 a_159_n91# a_n179_n179# a_63_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X3 a_n129_n91# a_n179_n179# a_n221_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_CBDHKH a_n33_n165# a_n189_n262# a_159_n165# a_n221_n165#
+ a_n129_n165# w_n263_n265# a_63_n165#
X0 a_n33_n165# a_n189_n262# a_n129_n165# w_n263_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X1 a_159_n165# a_n189_n262# a_63_n165# w_n263_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X2 a_63_n165# a_n189_n262# a_n33_n165# w_n263_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X3 a_n129_n165# a_n189_n262# a_n221_n165# w_n263_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_MRXJZU a_n321_n91# a_159_n91# a_351_n91# a_n33_n91#
+ a_n225_n91# a_n413_n91# a_63_n91# a_255_n91# a_n129_n91# a_n377_n179# VSUBS
X0 a_63_n91# a_n377_n179# a_n33_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X1 a_n33_n91# a_n377_n179# a_n129_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X2 a_351_n91# a_n377_n179# a_255_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X3 a_159_n91# a_n377_n179# a_63_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X4 a_255_n91# a_n377_n179# a_159_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X5 a_n321_n91# a_n377_n179# a_n413_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X6 a_n225_n91# a_n377_n179# a_n321_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X7 a_n129_n91# a_n377_n179# a_n225_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_CBVRKH a_n321_n165# a_n369_n262# a_n33_n165# w_n451_n265#
+ a_159_n165# a_255_n165# a_n413_n165# a_351_n165# a_n129_n165# a_63_n165# a_n225_n165#
X0 a_n33_n165# a_n369_n262# a_n129_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X1 a_351_n165# a_n369_n262# a_255_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X2 a_255_n165# a_n369_n262# a_159_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X3 a_n321_n165# a_n369_n262# a_n413_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X4 a_159_n165# a_n369_n262# a_63_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X5 a_n225_n165# a_n369_n262# a_n321_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X6 a_63_n165# a_n369_n262# a_n33_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X7 a_n129_n165# a_n369_n262# a_n225_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt capacitor_switch8 VDD Vin VSS Vout
XXM1 Vin VSS m1_90_960# VSS sky130_fd_pr__nfet_01v8_9CGS2F
XXM2 m1_90_960# Vin VDD VDD sky130_fd_pr__pfet_01v8_46WN3R
XXM3 VSS m1_90_960# m1_680_760# m1_680_760# VSS sky130_fd_pr__nfet_01v8_5XXJZ8
XXM4 VDD m1_680_760# VDD m1_680_760# m1_90_960# sky130_fd_pr__pfet_01v8_CBMBZG
XXM5 m1_1200_560# m1_1200_560# m1_1200_560# m1_680_760# VSS VSS VSS sky130_fd_pr__nfet_01v8_ZDVJZL
XXM6 m1_1200_560# m1_680_760# m1_1200_560# m1_1200_560# VDD VDD VDD sky130_fd_pr__pfet_01v8_CBDHKH
XXM7 VSS Vout Vout Vout Vout Vout VSS VSS VSS m1_1200_560# VSS sky130_fd_pr__nfet_01v8_MRXJZU
XXM8 VDD m1_1200_560# Vout VDD Vout VDD Vout Vout VDD VDD Vout sky130_fd_pr__pfet_01v8_CBVRKH
.ends

.subckt sky130_fd_sc_hd__diode_2 VGND VPWR DIODE VPB VNB
D0 VNB DIODE sky130_fd_pr__diode_pw2nd_05v5 pj=2.64e+06u area=4.347e+11p
.ends

.subckt sky130_fd_pr__nfet_01v8_ZZU2YL a_159_n91# a_n221_n91# a_n33_n91# a_n177_n179#
+ a_63_n91# a_n129_n91# VSUBS
X0 a_63_n91# a_n177_n179# a_n33_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X1 a_n33_n91# a_n177_n179# a_n129_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X2 a_159_n91# a_n177_n179# a_63_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X3 a_n129_n91# a_n177_n179# a_n221_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_C7DZJH a_n33_n165# a_n177_n262# w_n263_n295# a_159_n165#
+ a_n221_n165# a_n129_n165# a_63_n165#
X0 a_n33_n165# a_n177_n262# a_n129_n165# w_n263_n295# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X1 a_159_n165# a_n177_n262# a_63_n165# w_n263_n295# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X2 a_63_n165# a_n177_n262# a_n33_n165# w_n263_n295# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X3 a_n129_n165# a_n177_n262# a_n221_n165# w_n263_n295# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt capacitor_switch4 VDD Vin VSS Vout
Xsky130_fd_pr__pfet_01v8_46WN3R_0 m1_310_910# Vin VDD VDD sky130_fd_pr__pfet_01v8_46WN3R
Xsky130_fd_pr__nfet_01v8_ZZU2YL_0 VSS VSS VSS m1_310_910# Vout Vout VSS sky130_fd_pr__nfet_01v8_ZZU2YL
Xsky130_fd_pr__nfet_01v8_9CGS2F_0 Vin VSS m1_310_910# VSS sky130_fd_pr__nfet_01v8_9CGS2F
XXM4 VDD m1_310_910# VDD VDD VDD Vout Vout sky130_fd_pr__pfet_01v8_C7DZJH
.ends

.subckt sky130_fd_pr__pfet_01v8_S6MTYS a_n33_n165# w_n161_n265# a_n125_n165# a_63_n165#
+ a_n81_195#
X0 a_n33_n165# a_n81_195# a_n125_n165# w_n161_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X1 a_63_n165# a_n81_195# a_n33_n165# w_n161_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_9CME3F a_n73_n122# a_15_n122# a_n33_82# VSUBS
X0 a_15_n122# a_n33_82# a_n73_n122# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_Z2KCLS a_n33_173# a_n73_n213# a_15_n213# VSUBS
X0 a_15_n213# a_n33_173# a_n73_n213# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.82e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_5AWN3K a_15_n201# a_n33_160# a_n73_n201# w_n109_n263#
X0 a_15_n201# a_n33_160# a_n73_n201# w_n109_n263# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt capacitor_switch2 VDD Vin VSS Vout
Xsky130_fd_pr__pfet_01v8_S6MTYS_0 VDD VDD Vout Vout m1_n200_780# sky130_fd_pr__pfet_01v8_S6MTYS
XXM1 VSS m1_n200_780# Vin VSS sky130_fd_pr__nfet_01v8_9CME3F
XXM3 m1_n200_780# VSS Vout VSS sky130_fd_pr__nfet_01v8_Z2KCLS
Xsky130_fd_pr__pfet_01v8_5AWN3K_0 VDD Vin m1_n200_780# VDD sky130_fd_pr__pfet_01v8_5AWN3K
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_H9XL9H c1_n550_n500# m3_n650_n600#
X0 c1_n550_n500# m3_n650_n600# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
.ends

.subckt cap32 m4_4380_800# m4_5300_800# m4_5980_800# m4_500_800# m4_1180_800# m4_2100_800#
+ m4_2780_800# m4_3700_800#
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
.ends

.subckt cap8 m4_1180_800# m4_500_800#
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
.ends

.subckt cap64 m4_10100_800# m4_4380_800# m4_10780_800# m4_5300_800# m4_11700_800#
+ m4_5980_800# m4_500_800# m4_12380_800# m4_6900_800# m4_1180_800# m4_7580_800# m4_2100_800#
+ m4_8500_800# m4_2780_800# m4_9180_800# m4_3700_800#
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
.ends

.subckt cap4 m4_5300_0# m4_6000_0# m4_3700_0# m4_4400_0# m4_2100_0# m4_2800_0# m4_1200_0#
+ m4_500_0#
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0] m4_500_0# m4_1200_0# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1] m4_2100_0# m4_2800_0# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2] m4_3700_0# m4_4400_0# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3] m4_5300_0# m4_6000_0# sky130_fd_pr__cap_mim_m3_1_H9XL9H
.ends

.subckt cap16 m4_500_800# m4_1180_800# m4_2100_800# m4_2780_800#
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
.ends

.subckt cap2 m4_2100_0# m4_2800_0# m4_1200_0# m4_500_0#
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0] m4_500_0# m4_1200_0# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1] m4_2100_0# m4_2800_0# sky130_fd_pr__cap_mim_m3_1_H9XL9H
.ends

.subckt cap1 m4_1200_0# m4_500_0#
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0 m4_500_0# m4_1200_0# sky130_fd_pr__cap_mim_m3_1_H9XL9H
.ends

.subckt cap128 m4_10100_800# m4_17180_800# m4_16500_800# m4_23580_800# m4_22900_800#
+ m4_4380_800# m4_10780_800# m4_5300_800# m4_11700_800# m4_18780_800# m4_18100_800#
+ m4_24500_800# m4_25180_800# m4_5980_800# m4_500_800# m4_12380_800# m4_6900_800#
+ m4_13300_800# m4_20380_800# m4_19700_800# m4_1180_800# m4_7580_800# m4_2100_800#
+ m4_13980_800# m4_8500_800# m4_14900_800# m4_21980_800# m4_21300_800# m4_2780_800#
+ m4_9180_800# m4_3700_800# m4_15580_800#
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|0] m4_500_800# m4_1180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|1] m4_2100_800# m4_2780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|2] m4_3700_800# m4_4380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|3] m4_5300_800# m4_5980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|4] m4_6900_800# m4_7580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|5] m4_8500_800# m4_9180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|6] m4_10100_800# m4_10780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|7] m4_11700_800# m4_12380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|8] m4_13300_800# m4_13980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|8] m4_13300_800# m4_13980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|8] m4_13300_800# m4_13980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|8] m4_13300_800# m4_13980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|8] m4_13300_800# m4_13980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|8] m4_13300_800# m4_13980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|8] m4_13300_800# m4_13980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|8] m4_13300_800# m4_13980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|9] m4_14900_800# m4_15580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|9] m4_14900_800# m4_15580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|9] m4_14900_800# m4_15580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|9] m4_14900_800# m4_15580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|9] m4_14900_800# m4_15580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|9] m4_14900_800# m4_15580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|9] m4_14900_800# m4_15580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|9] m4_14900_800# m4_15580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|10] m4_16500_800# m4_17180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|10] m4_16500_800# m4_17180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|10] m4_16500_800# m4_17180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|10] m4_16500_800# m4_17180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|10] m4_16500_800# m4_17180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|10] m4_16500_800# m4_17180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|10] m4_16500_800# m4_17180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|10] m4_16500_800# m4_17180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|11] m4_18100_800# m4_18780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|11] m4_18100_800# m4_18780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|11] m4_18100_800# m4_18780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|11] m4_18100_800# m4_18780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|11] m4_18100_800# m4_18780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|11] m4_18100_800# m4_18780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|11] m4_18100_800# m4_18780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|11] m4_18100_800# m4_18780_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|12] m4_19700_800# m4_20380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|12] m4_19700_800# m4_20380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|12] m4_19700_800# m4_20380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|12] m4_19700_800# m4_20380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|12] m4_19700_800# m4_20380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|12] m4_19700_800# m4_20380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|12] m4_19700_800# m4_20380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|12] m4_19700_800# m4_20380_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|13] m4_21300_800# m4_21980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|13] m4_21300_800# m4_21980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|13] m4_21300_800# m4_21980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|13] m4_21300_800# m4_21980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|13] m4_21300_800# m4_21980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|13] m4_21300_800# m4_21980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|13] m4_21300_800# m4_21980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|13] m4_21300_800# m4_21980_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|14] m4_22900_800# m4_23580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|14] m4_22900_800# m4_23580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|14] m4_22900_800# m4_23580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|14] m4_22900_800# m4_23580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|14] m4_22900_800# m4_23580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|14] m4_22900_800# m4_23580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|14] m4_22900_800# m4_23580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|14] m4_22900_800# m4_23580_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[0|15] m4_24500_800# m4_25180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[1|15] m4_24500_800# m4_25180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[2|15] m4_24500_800# m4_25180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[3|15] m4_24500_800# m4_25180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[4|15] m4_24500_800# m4_25180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[5|15] m4_24500_800# m4_25180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[6|15] m4_24500_800# m4_25180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
Xsky130_fd_pr__cap_mim_m3_1_H9XL9H_0[7|15] m4_24500_800# m4_25180_800# sky130_fd_pr__cap_mim_m3_1_H9XL9H
.ends

.subckt capacitor_array sw_sp_n9 sw_sp_n8 sw_sp_n7 sw_sp_n6 sw_sp_n5 sw_sp_n4 sw_sp_n3
+ sw_sp_n2 sw_sp_n1 Vin_p Vin_n sw_sp_p9 sw_sp_p8 sw_sp_p7 sw_sp_p6 sw_sp_p5 sw_sp_p4
+ sw_sp_p3 sw_sp_p2 sw_sp_p1 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3 sw_p2 sw_p1 sw_n8
+ sw_n7 sw_n6 sw_n5 sw_n4 sw_n3 sw_n2 sw_n1
Xcap32_1 Vin_p sw_p3 Vin_p sw_p3 Vin_p sw_p3 Vin_p sw_p3 cap32
Xcap8_3 Vin_n sw_sp_n5 cap8
Xcap64_3 sw_sp_n2 Vin_n Vin_n sw_sp_n2 sw_sp_n2 Vin_n sw_sp_n2 Vin_n sw_sp_n2 Vin_n
+ Vin_n sw_sp_n2 sw_sp_n2 Vin_n Vin_n sw_sp_n2 cap64
Xcap32_2 Vin_n sw_n3 Vin_n sw_n3 Vin_n sw_n3 Vin_n sw_n3 cap32
Xcap32_3 Vin_n sw_sp_n3 Vin_n sw_sp_n3 Vin_n sw_sp_n3 Vin_n sw_sp_n3 cap32
Xcap4_0 sw_sp_p6 Vin_p sw_sp_p6 Vin_p sw_sp_p6 Vin_p Vin_p sw_sp_p6 cap4
Xcap4_1 sw_p6 Vin_p sw_p6 Vin_p sw_p6 Vin_p Vin_p sw_p6 cap4
Xcap16_0 sw_sp_p4 Vin_p sw_sp_p4 Vin_p cap16
Xcap16_1 sw_p4 Vin_p sw_p4 Vin_p cap16
Xcap4_2 sw_n6 Vin_n sw_n6 Vin_n sw_n6 Vin_n Vin_n sw_n6 cap4
Xcap16_2 sw_n4 Vin_n sw_n4 Vin_n cap16
Xcap2_0 sw_sp_p7 Vin_p Vin_p sw_sp_p7 cap2
Xcap4_3 sw_sp_n6 Vin_n sw_sp_n6 Vin_n sw_sp_n6 Vin_n Vin_n sw_sp_n6 cap4
Xcap16_3 sw_sp_n4 Vin_n sw_sp_n4 Vin_n cap16
Xcap2_1 sw_n7 Vin_n Vin_n sw_n7 cap2
Xcap2_2 sw_sp_n7 Vin_n Vin_n sw_sp_n7 cap2
Xcap2_3 sw_p7 Vin_p Vin_p sw_p7 cap2
Xcap1_0 Vin_p sw_sp_p8 cap1
Xcap1_1 Vin_n sw_n8 cap1
Xcap1_2 Vin_n sw_sp_n9 cap1
Xcap128_0 sw_sp_p1 Vin_p sw_sp_p1 Vin_p sw_sp_p1 Vin_p Vin_p sw_sp_p1 sw_sp_p1 Vin_p
+ sw_sp_p1 sw_sp_p1 Vin_p Vin_p sw_sp_p1 Vin_p sw_sp_p1 sw_sp_p1 Vin_p sw_sp_p1 Vin_p
+ Vin_p sw_sp_p1 Vin_p sw_sp_p1 sw_sp_p1 Vin_p sw_sp_p1 Vin_p Vin_p sw_sp_p1 Vin_p
+ cap128
Xcap1_3 Vin_n sw_sp_n8 cap1
Xcap1_4 Vin_p sw_sp_p9 cap1
Xcap128_1 sw_p1 Vin_p sw_p1 Vin_p sw_p1 Vin_p Vin_p sw_p1 sw_p1 Vin_p sw_p1 sw_p1
+ Vin_p Vin_p sw_p1 Vin_p sw_p1 sw_p1 Vin_p sw_p1 Vin_p Vin_p sw_p1 Vin_p sw_p1 sw_p1
+ Vin_p sw_p1 Vin_p Vin_p sw_p1 Vin_p cap128
Xcap128_2 sw_n1 Vin_n sw_n1 Vin_n sw_n1 Vin_n Vin_n sw_n1 sw_n1 Vin_n sw_n1 sw_n1
+ Vin_n Vin_n sw_n1 Vin_n sw_n1 sw_n1 Vin_n sw_n1 Vin_n Vin_n sw_n1 Vin_n sw_n1 sw_n1
+ Vin_n sw_n1 Vin_n Vin_n sw_n1 Vin_n cap128
Xcap1_5 Vin_p sw_p8 cap1
Xcap128_3 sw_sp_n1 Vin_n sw_sp_n1 Vin_n sw_sp_n1 Vin_n Vin_n sw_sp_n1 sw_sp_n1 Vin_n
+ sw_sp_n1 sw_sp_n1 Vin_n Vin_n sw_sp_n1 Vin_n sw_sp_n1 sw_sp_n1 Vin_n sw_sp_n1 Vin_n
+ Vin_n sw_sp_n1 Vin_n sw_sp_n1 sw_sp_n1 Vin_n sw_sp_n1 Vin_n Vin_n sw_sp_n1 Vin_n
+ cap128
Xcap64_0 sw_p2 Vin_p Vin_p sw_p2 sw_p2 Vin_p sw_p2 Vin_p sw_p2 Vin_p Vin_p sw_p2 sw_p2
+ Vin_p Vin_p sw_p2 cap64
Xcap8_0 Vin_p sw_sp_p5 cap8
Xcap64_1 sw_sp_p2 Vin_p Vin_p sw_sp_p2 sw_sp_p2 Vin_p sw_sp_p2 Vin_p sw_sp_p2 Vin_p
+ Vin_p sw_sp_p2 sw_sp_p2 Vin_p Vin_p sw_sp_p2 cap64
Xcap8_1 Vin_p sw_p5 cap8
Xcap32_0 Vin_p sw_sp_p3 Vin_p sw_sp_p3 Vin_p sw_sp_p3 Vin_p sw_sp_p3 cap32
Xcap8_2 Vin_n sw_n5 cap8
Xcap64_2 sw_n2 Vin_n Vin_n sw_n2 sw_n2 Vin_n sw_n2 Vin_n sw_n2 Vin_n Vin_n sw_n2 sw_n2
+ Vin_n Vin_n sw_n2 cap64
.ends

.subckt sky130_fd_sc_hd__bufbuf_16 VGND VPWR A X VNB VPB
X0 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_109_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 a_549_47# a_215_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X21 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X31 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 VGND a_215_47# a_549_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X34 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X35 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 VGND a_549_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 a_215_47# a_109_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X40 a_215_47# a_109_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X41 VPWR a_109_47# a_215_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X42 X a_549_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 VPWR a_215_47# a_549_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X45 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X46 a_109_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_549_47# a_215_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 VPWR a_549_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_109_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X51 X a_549_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_BBAHKR a_n33_n165# a_159_n165# a_n179_n262# a_n221_n165#
+ a_n129_n165# w_n263_n265# a_63_n165#
X0 a_n33_n165# a_n179_n262# a_n129_n165# w_n263_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X1 a_159_n165# a_n179_n262# a_63_n165# w_n263_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X2 a_63_n165# a_n179_n262# a_n33_n165# w_n263_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X3 a_n129_n165# a_n179_n262# a_n221_n165# w_n263_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_HRFJZU a_n321_n91# a_n369_n179# a_159_n91# a_351_n91#
+ a_n33_n91# a_n225_n91# a_n413_n91# a_63_n91# a_255_n91# a_n129_n91# VSUBS
X0 a_63_n91# a_n369_n179# a_n33_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X1 a_n33_n91# a_n369_n179# a_n129_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X2 a_351_n91# a_n369_n179# a_255_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X3 a_159_n91# a_n369_n179# a_63_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X4 a_255_n91# a_n369_n179# a_159_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X5 a_n321_n91# a_n369_n179# a_n413_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X6 a_n225_n91# a_n369_n179# a_n321_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X7 a_n129_n91# a_n369_n179# a_n225_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_5EDJZL a_159_n91# a_n221_n91# a_n33_n91# a_n179_n179#
+ a_63_n91# a_n129_n91# VSUBS
X0 a_63_n91# a_n179_n179# a_n33_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X1 a_n33_n91# a_n179_n179# a_n129_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X2 a_159_n91# a_n179_n179# a_63_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X3 a_n129_n91# a_n179_n179# a_n221_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_BBSRKR a_n321_n165# a_n33_n165# w_n451_n265# a_159_n165#
+ a_255_n165# a_n413_n165# a_351_n165# a_n129_n165# a_63_n165# a_n225_n165# a_n377_n262#
X0 a_n33_n165# a_n377_n262# a_n129_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X1 a_351_n165# a_n377_n262# a_255_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X2 a_255_n165# a_n377_n262# a_159_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X3 a_n321_n165# a_n377_n262# a_n413_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X4 a_159_n165# a_n377_n262# a_63_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X5 a_n225_n165# a_n377_n262# a_n321_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X6 a_63_n165# a_n377_n262# a_n33_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X7 a_n129_n165# a_n377_n262# a_n225_n165# w_n451_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_29RM5N a_n609_n91# a_447_n91# a_n321_n91# a_n753_n179#
+ a_159_n91# a_639_n91# a_n513_n91# a_351_n91# a_n33_n91# a_n797_n91# a_n225_n91#
+ a_n705_n91# a_543_n91# a_63_n91# a_n417_n91# a_255_n91# a_735_n91# a_n129_n91# VSUBS
X0 a_n609_n91# a_n753_n179# a_n705_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X1 a_63_n91# a_n753_n179# a_n33_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X2 a_n33_n91# a_n753_n179# a_n129_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X3 a_351_n91# a_n753_n179# a_255_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X4 a_159_n91# a_n753_n179# a_63_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X5 a_255_n91# a_n753_n179# a_159_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X6 a_447_n91# a_n753_n179# a_351_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X7 a_543_n91# a_n753_n179# a_447_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X8 a_735_n91# a_n753_n179# a_639_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X9 a_639_n91# a_n753_n179# a_543_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X10 a_n321_n91# a_n753_n179# a_n417_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X11 a_n705_n91# a_n753_n179# a_n797_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X12 a_n513_n91# a_n753_n179# a_n609_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X13 a_n417_n91# a_n753_n179# a_n513_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X14 a_n225_n91# a_n753_n179# a_n321_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X15 a_n129_n91# a_n753_n179# a_n225_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_2FR7QD a_n321_n165# a_639_n165# a_n753_n262# a_735_n165#
+ a_n33_n165# a_447_n165# a_543_n165# a_159_n165# a_n609_n165# a_255_n165# a_n705_n165#
+ a_351_n165# a_n417_n165# a_n129_n165# a_n513_n165# a_63_n165# a_n225_n165# a_n797_n165#
+ w_n837_n265#
X0 a_639_n165# a_n753_n262# a_543_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X1 a_n705_n165# a_n753_n262# a_n797_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X2 a_n33_n165# a_n753_n262# a_n129_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X3 a_351_n165# a_n753_n262# a_255_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X4 a_n609_n165# a_n753_n262# a_n705_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X5 a_255_n165# a_n753_n262# a_159_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X6 a_n321_n165# a_n753_n262# a_n417_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X7 a_543_n165# a_n753_n262# a_447_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X8 a_159_n165# a_n753_n262# a_63_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X9 a_n225_n165# a_n753_n262# a_n321_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X10 a_447_n165# a_n753_n262# a_351_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X11 a_n513_n165# a_n753_n262# a_n609_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X12 a_63_n165# a_n753_n262# a_n33_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X13 a_735_n165# a_n753_n262# a_639_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X14 a_n129_n165# a_n753_n262# a_n225_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
X15 a_n417_n165# a_n753_n262# a_n513_n165# w_n837_n265# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.65e+06u l=150000u
.ends

.subckt capacitor_switch16 VDD Vin VSS Vout
Xsky130_fd_pr__pfet_01v8_46WN3R_0 m1_n190_980# Vin VDD VDD sky130_fd_pr__pfet_01v8_46WN3R
Xsky130_fd_pr__nfet_01v8_9CGS2F_0 Vin VSS m1_n190_980# VSS sky130_fd_pr__nfet_01v8_9CGS2F
XXM4 m1_430_590# m1_430_590# m1_n190_980# m1_430_590# VDD VDD VDD sky130_fd_pr__pfet_01v8_BBAHKR
XXM5 VSS m1_430_590# m1_930_200# m1_930_200# m1_930_200# m1_930_200# m1_930_200# VSS
+ VSS VSS VSS sky130_fd_pr__nfet_01v8_HRFJZU
Xsky130_fd_pr__nfet_01v8_5EDJZL_0 m1_430_590# m1_430_590# m1_430_590# m1_n190_980#
+ VSS VSS VSS sky130_fd_pr__nfet_01v8_5EDJZL
XXM6 VDD m1_930_200# VDD m1_930_200# VDD m1_930_200# m1_930_200# VDD VDD m1_930_200#
+ m1_430_590# sky130_fd_pr__pfet_01v8_BBSRKR
XXM7 Vout VSS VSS m1_930_200# Vout VSS VSS Vout Vout Vout Vout VSS Vout VSS Vout VSS
+ Vout VSS VSS sky130_fd_pr__nfet_01v8_29RM5N
XXM8 VDD VDD m1_930_200# Vout Vout VDD Vout Vout Vout VDD VDD Vout Vout VDD VDD VDD
+ Vout Vout VDD sky130_fd_pr__pfet_01v8_2FR7QD
.ends

.subckt dac sw_sp_n9 sw_sp_n8 sw_sp_n7 sw_sp_n6 sw_sp_n5 sw_sp_n4 sw_sp_n3 sw_sp_n2
+ sw_sp_n1 sw_sp_p9 sw_sp_p8 sw_sp_p7 sw_sp_p6 sw_sp_p5 sw_sp_p4 sw_sp_p3 sw_sp_p2
+ sw_sp_p1 sw_n8 sw_n7 sw_n6 sw_n5 sw_n4 sw_n3 sw_n2 sw_n1 sw_p8 sw_p7 sw_p6 sw_p5
+ sw_p4 sw_p3 sw_p2 sw_p1 sample_sw_buf_in sample_sw_buf_out VDD Vin_p Vin_n VSS
Xcapacitor_switch8_7 VDD capacitor_switch8_7/Vin VSS capacitor_array_0/sw_p4 capacitor_switch8
Xsky130_fd_sc_hd__diode_2_34 VSS VDD capacitor_switch8_6/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_12 VSS VDD capacitor_switch8_2/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch4_1 VDD sw_n6 VSS capacitor_array_0/sw_n6 capacitor_switch4
Xsky130_fd_sc_hd__diode_2_23 VSS VDD sw_p2 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_35 VSS VDD capacitor_switch4_7/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch4_2 VDD capacitor_switch4_2/Vin VSS capacitor_switch4_2/Vout capacitor_switch4
Xsky130_fd_sc_hd__diode_2_13 VSS VDD capacitor_switch8_3/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_24 VSS VDD sw_sp_p4 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_36 VSS VDD capacitor_switch16_5/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_14 VSS VDD capacitor_switch4_0/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_25 VSS VDD sw_sp_p2 VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch4_3 VDD sw_sp_n6 VSS capacitor_switch4_3/Vout capacitor_switch4
Xcapacitor_switch2_0 VDD sw_sp_n9 VSS capacitor_switch2_0/Vout capacitor_switch2
Xsky130_fd_sc_hd__diode_2_37 VSS VDD capacitor_switch8_5/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_15 VSS VDD capacitor_switch16_2/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch4_4 VDD sw_sp_p6 VSS capacitor_switch4_4/Vout capacitor_switch4
Xsky130_fd_sc_hd__diode_2_26 VSS VDD sw_p4 VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch2_1 VDD sw_sp_n7 VSS capacitor_switch2_1/Vout capacitor_switch2
Xsky130_fd_sc_hd__diode_2_38 VSS VDD capacitor_switch16_3/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_16 VSS VDD capacitor_switch16_1/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_27 VSS VDD sw_sp_p5 VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch2_2 VDD sw_sp_n8 VSS capacitor_switch2_2/Vout capacitor_switch2
Xcapacitor_switch4_5 VDD sw_p6 VSS capacitor_array_0/sw_p6 capacitor_switch4
Xsky130_fd_sc_hd__diode_2_39 VSS VDD capacitor_switch16_6/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch4_6 VDD capacitor_switch4_6/Vin VSS capacitor_array_0/sw_p5 capacitor_switch4
Xsky130_fd_sc_hd__diode_2_17 VSS VDD capacitor_switch16_7/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_28 VSS VDD sw_sp_p3 VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch2_3 VDD sw_n7 VSS capacitor_array_0/sw_n7 capacitor_switch2
Xsky130_fd_sc_hd__diode_2_18 VSS VDD capacitor_switch16_0/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_29 VSS VDD sample_sw_buf_in VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch2_4 VDD sw_n8 VSS capacitor_array_0/sw_n8 capacitor_switch2
Xcapacitor_switch4_7 VDD capacitor_switch4_7/Vin VSS capacitor_switch4_7/Vout capacitor_switch4
Xsky130_fd_sc_hd__diode_2_19 VSS VDD capacitor_switch8_1/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch2_5 VDD sw_sp_p8 VSS capacitor_switch2_5/Vout capacitor_switch2
Xcapacitor_array_0 capacitor_switch2_0/Vout capacitor_switch2_2/Vout capacitor_switch2_1/Vout
+ capacitor_switch4_3/Vout capacitor_switch4_2/Vout capacitor_switch8_0/Vout capacitor_switch8_1/Vout
+ capacitor_switch16_1/Vout capacitor_switch16_2/Vout Vin_p Vin_n capacitor_switch2_9/Vout
+ capacitor_switch2_5/Vout capacitor_switch2_6/Vout capacitor_switch4_4/Vout capacitor_switch4_7/Vout
+ capacitor_switch8_6/Vout capacitor_switch8_5/Vout capacitor_switch16_3/Vout capacitor_switch16_4/Vout
+ capacitor_array_0/sw_p8 capacitor_array_0/sw_p7 capacitor_array_0/sw_p6 capacitor_array_0/sw_p5
+ capacitor_array_0/sw_p4 capacitor_array_0/sw_p3 capacitor_array_0/sw_p2 capacitor_array_0/sw_p1
+ capacitor_array_0/sw_n8 capacitor_array_0/sw_n7 capacitor_array_0/sw_n6 capacitor_array_0/sw_n5
+ capacitor_array_0/sw_n4 capacitor_array_0/sw_n3 capacitor_array_0/sw_n2 capacitor_array_0/sw_n1
+ capacitor_array
Xcapacitor_switch2_6 VDD sw_sp_p7 VSS capacitor_switch2_6/Vout capacitor_switch2
Xcapacitor_switch2_7 VDD sw_p7 VSS capacitor_array_0/sw_p7 capacitor_switch2
Xcapacitor_switch2_8 VDD sw_p8 VSS capacitor_array_0/sw_p8 capacitor_switch2
Xcapacitor_switch2_9 VDD sw_sp_p9 VSS capacitor_switch2_9/Vout capacitor_switch2
Xsky130_fd_sc_hd__bufbuf_16_20 VSS VDD sw_sp_p2 capacitor_switch16_3/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_21 VSS VDD sample_sw_buf_in sky130_fd_sc_hd__bufbuf_16_21/X
+ VSS VDD sky130_fd_sc_hd__bufbuf_16
Xcapacitor_switch16_0 VDD capacitor_switch16_0/Vin VSS capacitor_array_0/sw_n2 capacitor_switch16
Xsky130_fd_sc_hd__bufbuf_16_0 VSS VDD sw_n4 capacitor_switch8_3/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_10 VSS VDD sky130_fd_sc_hd__bufbuf_16_21/X sample_sw_buf_out
+ VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_11 VSS VDD sw_p4 capacitor_switch8_7/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xcapacitor_switch16_1 VDD capacitor_switch16_1/Vin VSS capacitor_switch16_1/Vout capacitor_switch16
Xsky130_fd_sc_hd__bufbuf_16_1 VSS VDD sw_n2 capacitor_switch16_0/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_12 VSS VDD sw_p3 capacitor_switch8_4/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xcapacitor_switch16_2 VDD capacitor_switch16_2/Vin VSS capacitor_switch16_2/Vout capacitor_switch16
Xsky130_fd_sc_hd__bufbuf_16_2 VSS VDD sw_sp_n4 capacitor_switch8_0/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_13 VSS VDD sw_p5 capacitor_switch4_6/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_3 VSS VDD sw_n3 capacitor_switch8_2/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xcapacitor_switch16_3 VDD capacitor_switch16_3/Vin VSS capacitor_switch16_3/Vout capacitor_switch16
Xsky130_fd_sc_hd__bufbuf_16_14 VSS VDD sw_sp_p5 capacitor_switch4_7/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_4 VSS VDD sw_n5 capacitor_switch4_0/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xcapacitor_switch16_4 VDD capacitor_switch16_4/Vin VSS capacitor_switch16_4/Vout capacitor_switch16
Xsky130_fd_sc_hd__bufbuf_16_15 VSS VDD sw_sp_p4 capacitor_switch8_6/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_5 VSS VDD sw_sp_n1 capacitor_switch16_2/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xcapacitor_switch16_5 VDD capacitor_switch16_5/Vin VSS capacitor_array_0/sw_p2 capacitor_switch16
Xsky130_fd_sc_hd__diode_2_0 VSS VDD sw_sp_n1 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__bufbuf_16_16 VSS VDD sw_sp_p3 capacitor_switch8_5/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_6 VSS VDD sw_sp_n3 capacitor_switch8_1/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xcapacitor_switch16_6 VDD capacitor_switch16_6/Vin VSS capacitor_array_0/sw_p1 capacitor_switch16
Xsky130_fd_sc_hd__diode_2_1 VSS VDD sw_sp_n2 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__bufbuf_16_17 VSS VDD sw_p2 capacitor_switch16_5/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xcapacitor_switch16_7 VDD capacitor_switch16_7/Vin VSS capacitor_array_0/sw_n1 capacitor_switch16
Xsky130_fd_sc_hd__bufbuf_16_7 VSS VDD sw_sp_n5 capacitor_switch4_2/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__diode_2_2 VSS VDD sw_n1 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__bufbuf_16_18 VSS VDD sw_sp_p1 capacitor_switch16_4/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_8 VSS VDD sw_n1 capacitor_switch16_7/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__diode_2_3 VSS VDD sw_n2 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__bufbuf_16_19 VSS VDD sw_p1 capacitor_switch16_6/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__bufbuf_16_9 VSS VDD sw_sp_n2 capacitor_switch16_1/Vin VSS VDD sky130_fd_sc_hd__bufbuf_16
Xsky130_fd_sc_hd__diode_2_4 VSS VDD sw_sp_n3 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_5 VSS VDD sw_sp_n4 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_6 VSS VDD sw_sp_n5 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_7 VSS VDD sw_n3 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_8 VSS VDD sw_n5 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_9 VSS VDD sw_n4 VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch8_0 VDD capacitor_switch8_0/Vin VSS capacitor_switch8_0/Vout capacitor_switch8
Xcapacitor_switch8_1 VDD capacitor_switch8_1/Vin VSS capacitor_switch8_1/Vout capacitor_switch8
Xcapacitor_switch8_2 VDD capacitor_switch8_2/Vin VSS capacitor_array_0/sw_n3 capacitor_switch8
Xsky130_fd_sc_hd__diode_2_40 VSS VDD capacitor_switch16_4/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch8_3 VDD capacitor_switch8_3/Vin VSS capacitor_array_0/sw_n4 capacitor_switch8
Xsky130_fd_sc_hd__diode_2_30 VSS VDD sw_p1 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_41 VSS VDD sw_sp_p1 VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch8_4 VDD capacitor_switch8_4/Vin VSS capacitor_array_0/sw_p3 capacitor_switch8
Xsky130_fd_sc_hd__diode_2_42 VSS VDD sky130_fd_sc_hd__bufbuf_16_21/X VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_31 VSS VDD capacitor_switch4_6/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_20 VSS VDD sample_sw_buf_out VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch8_5 VDD capacitor_switch8_5/Vin VSS capacitor_switch8_5/Vout capacitor_switch8
Xsky130_fd_sc_hd__diode_2_32 VSS VDD capacitor_switch8_4/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_10 VSS VDD capacitor_switch8_0/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_21 VSS VDD sw_p3 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_33 VSS VDD capacitor_switch8_7/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_11 VSS VDD capacitor_switch4_2/Vin VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_22 VSS VDD sw_p5 VDD VSS sky130_fd_sc_hd__diode_2
Xcapacitor_switch8_6 VDD capacitor_switch8_6/Vin VSS capacitor_switch8_6/Vout capacitor_switch8
Xcapacitor_switch4_0 VDD capacitor_switch4_0/Vin VSS capacitor_array_0/sw_n5 capacitor_switch4
.ends

.subckt sky130_fd_pr__nfet_01v8_MRUJZ4 a_n321_n91# a_159_n91# a_351_n91# a_n33_n91#
+ a_n225_n91# a_n413_n91# a_63_n91# a_255_n91# a_n129_n91# a_n377_n179# VSUBS
X0 a_63_n91# a_n377_n179# a_n33_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X1 a_n33_n91# a_n377_n179# a_n129_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X2 a_351_n91# a_n377_n179# a_255_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X3 a_159_n91# a_n377_n179# a_63_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X4 a_255_n91# a_n377_n179# a_159_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X5 a_n321_n91# a_n377_n179# a_n413_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X6 a_n225_n91# a_n377_n179# a_n321_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X7 a_n129_n91# a_n377_n179# a_n225_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_6ZNTNB c1_n1050_n1000# m3_n1150_n1100#
X0 c1_n1050_n1000# m3_n1150_n1100# sky130_fd_pr__cap_mim_m3_1 l=1e+07u w=1e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_E9NJWS a_n73_n125# a_n33_n222# a_15_n125# w_n109_n225#
X0 a_15_n125# a_n33_n222# a_n73_n125# w_n109_n225# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_SKSN8V a_n73_n197# a_n33_156# w_n109_n259# a_15_n197#
X0 a_15_n197# a_n33_156# a_n73_n197# w_n109_n259# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ZWFJZ8 a_n33_n91# a_63_n91# a_n125_n91# a_n85_n179#
+ VSUBS
X0 a_63_n91# a_n85_n179# a_n33_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
X1 a_n33_n91# a_n85_n179# a_n125_n91# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=910000u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_P7BBP7 a_n369_n455# a_303_n455# a_n465_n455# a_n708_n543#
+ a_15_n455# a_n561_n455# a_n177_n455# a_111_n455# a_n273_n455# a_n749_n455# a_687_n455#
+ a_399_n455# a_n81_n455# a_495_n455# a_591_n455# a_n657_n455# a_207_n455# VSUBS
X0 a_n273_n455# a_n708_n543# a_n369_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X1 a_591_n455# a_n708_n543# a_495_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X2 a_207_n455# a_n708_n543# a_111_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X3 a_n177_n455# a_n708_n543# a_n273_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X4 a_495_n455# a_n708_n543# a_399_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X5 a_n561_n455# a_n708_n543# a_n657_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X6 a_111_n455# a_n708_n543# a_15_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X7 a_399_n455# a_n708_n543# a_303_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X8 a_n465_n455# a_n708_n543# a_n561_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X9 a_687_n455# a_n708_n543# a_591_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X10 a_n81_n455# a_n708_n543# a_n177_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X11 a_15_n455# a_n708_n543# a_n81_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X12 a_n369_n455# a_n708_n543# a_n465_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X13 a_n657_n455# a_n708_n543# a_n749_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
X14 a_303_n455# a_n708_n543# a_207_n455# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.55e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_RQ978N a_207_n100# a_15_n100# a_n177_n100# a_111_n100#
+ a_n225_n197# w_n305_n200# a_n81_n100# a_n269_n100#
X0 a_207_n100# a_n225_n197# a_111_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_15_n100# a_n225_n197# a_n81_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_111_n100# a_n225_n197# a_15_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_n81_n100# a_n225_n197# a_n177_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_n177_n100# a_n225_n197# a_n269_n100# w_n305_n200# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt bootstrapped_sampling_switch Vin_p Vin_n VDD VSS Clk Vout_n Vout_p
Xsky130_fd_pr__nfet_01v8_9CME3F_0 m1_4790_n3480# m1_4820_n4010# m1_5270_n4710# VSS
+ sky130_fd_pr__nfet_01v8_9CME3F
Xsky130_fd_pr__nfet_01v8_9CME3F_2 m1_7920_n3050# VSS m1_7860_n2950# VSS sky130_fd_pr__nfet_01v8_9CME3F
Xsky130_fd_pr__nfet_01v8_9CME3F_1 m1_5360_n3070# VSS m1_4560_n3710# VSS sky130_fd_pr__nfet_01v8_9CME3F
Xsky130_fd_pr__nfet_01v8_9CME3F_3 m1_8270_n4840# m1_8070_n5070# m1_7900_n4710# VSS
+ sky130_fd_pr__nfet_01v8_9CME3F
Xsky130_fd_pr__nfet_01v8_MRUJZ4_0 VSS m1_8070_n5070# m1_8070_n5070# m1_8070_n5070#
+ m1_8070_n5070# m1_8070_n5070# VSS VSS VSS m1_7860_n2950# VSS sky130_fd_pr__nfet_01v8_MRUJZ4
Xsky130_fd_pr__nfet_01v8_9CGS2F_0 m1_5270_n4710# m1_4820_n4010# Vin_n VSS sky130_fd_pr__nfet_01v8_9CGS2F
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_0[0|0] m1_4820_n4010# w_5020_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_0[1|0] m1_4820_n4010# w_5020_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_0[2|0] m1_4820_n4010# w_5020_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_0[0|1] m1_4820_n4010# w_5020_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_0[1|1] m1_4820_n4010# w_5020_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_0[2|1] m1_4820_n4010# w_5020_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_0[0|2] m1_4820_n4010# w_5020_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_0[1|2] m1_4820_n4010# w_5020_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_0[2|2] m1_4820_n4010# w_5020_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_1[0|0] m1_8070_n5070# w_8000_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_1[1|0] m1_8070_n5070# w_8000_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_1[2|0] m1_8070_n5070# w_8000_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_1[0|1] m1_8070_n5070# w_8000_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_1[1|1] m1_8070_n5070# w_8000_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_1[2|1] m1_8070_n5070# w_8000_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_1[0|2] m1_8070_n5070# w_8000_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_1[1|2] m1_8070_n5070# w_8000_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__cap_mim_m3_1_6ZNTNB_1[2|2] m1_8070_n5070# w_8000_n4620# sky130_fd_pr__cap_mim_m3_1_6ZNTNB
Xsky130_fd_pr__nfet_01v8_9CGS2F_2 Clk m1_4560_n3710# VSS VSS sky130_fd_pr__nfet_01v8_9CGS2F
Xsky130_fd_pr__nfet_01v8_9CGS2F_1 Clk m1_4820_n4010# m1_4790_n3480# VSS sky130_fd_pr__nfet_01v8_9CGS2F
Xsky130_fd_pr__nfet_01v8_9CGS2F_3 Clk m1_7860_n2950# VSS VSS sky130_fd_pr__nfet_01v8_9CGS2F
XXM1 VSS m1_4820_n4010# m1_4820_n4010# m1_4820_n4010# m1_4820_n4010# m1_4820_n4010#
+ VSS VSS VSS m1_4560_n3710# VSS sky130_fd_pr__nfet_01v8_MRUJZ4
XXM2 m1_4790_n3480# Clk VDD VDD sky130_fd_pr__pfet_01v8_E9NJWS
Xsky130_fd_pr__nfet_01v8_9CGS2F_4 m1_7900_n4710# m1_8070_n5070# Vin_p VSS sky130_fd_pr__nfet_01v8_9CGS2F
Xsky130_fd_pr__nfet_01v8_9CGS2F_5 Clk m1_8070_n5070# m1_8270_n4840# VSS sky130_fd_pr__nfet_01v8_9CGS2F
XXM5 m1_5270_n4710# m1_4790_n3480# w_5020_n4620# w_5020_n4620# sky130_fd_pr__pfet_01v8_SKSN8V
XXM9 m1_5360_n3070# m1_5270_n4710# m1_5270_n4710# VDD VSS sky130_fd_pr__nfet_01v8_ZWFJZ8
XXM8 Vin_n Vout_n Vout_n m1_5270_n4710# Vin_n Vin_n Vin_n Vout_n Vout_n Vin_n Vout_n
+ Vin_n Vout_n Vout_n Vin_n Vout_n Vin_n VSS sky130_fd_pr__nfet_01v8_P7BBP7
Xsky130_fd_pr__pfet_01v8_SKSN8V_0 m1_7900_n4710# m1_8270_n4840# w_8000_n4620# w_8000_n4620#
+ sky130_fd_pr__pfet_01v8_SKSN8V
Xsky130_fd_pr__pfet_01v8_RQ978N_0 w_5020_n4620# w_5020_n4620# w_5020_n4620# VDD m1_5270_n4710#
+ w_5020_n4620# VDD VDD sky130_fd_pr__pfet_01v8_RQ978N
Xsky130_fd_pr__pfet_01v8_E9NJWS_0 m1_4560_n3710# Clk VDD VDD sky130_fd_pr__pfet_01v8_E9NJWS
Xsky130_fd_pr__pfet_01v8_RQ978N_1 w_8000_n4620# w_8000_n4620# w_8000_n4620# VDD m1_7900_n4710#
+ w_8000_n4620# VDD VDD sky130_fd_pr__pfet_01v8_RQ978N
Xsky130_fd_pr__pfet_01v8_E9NJWS_1 m1_7860_n2950# Clk VDD VDD sky130_fd_pr__pfet_01v8_E9NJWS
Xsky130_fd_pr__pfet_01v8_E9NJWS_2 m1_8270_n4840# Clk VDD VDD sky130_fd_pr__pfet_01v8_E9NJWS
Xsky130_fd_pr__nfet_01v8_ZWFJZ8_0 m1_7920_n3050# m1_7900_n4710# m1_7900_n4710# VDD
+ VSS sky130_fd_pr__nfet_01v8_ZWFJZ8
Xsky130_fd_pr__nfet_01v8_P7BBP7_0 Vin_p Vout_p Vout_p m1_7900_n4710# Vin_p Vin_p Vin_p
+ Vout_p Vout_p Vin_p Vout_p Vin_p Vout_p Vout_p Vin_p Vout_p Vin_p VSS sky130_fd_pr__nfet_01v8_P7BBP7
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_8 VGND VPWR A X VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkdlybuf4s15_1 VGND VPWR A X VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_282_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_394_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_282_47# a_394_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 X a_394_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_282_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=150000u
X6 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_282_47# a_394_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=820000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_QPTUVJ a_n33_n161# a_159_n161# a_n191_n258# w_n257_n271#
+ a_n221_n161# a_n129_n161# a_63_n161#
X0 a_159_n161# a_n191_n258# a_63_n161# w_n257_n271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X1 a_63_n161# a_n191_n258# a_n33_n161# w_n257_n271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X2 a_n129_n161# a_n191_n258# a_n221_n161# w_n257_n271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X3 a_n33_n161# a_n191_n258# a_n129_n161# w_n257_n271# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_FBQ47L a_63_n500# a_n33_n500# a_n81_n597# w_n161_n600#
+ a_n125_n500#
X0 a_n33_n500# a_n81_n597# a_n125_n500# w_n161_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1 a_63_n500# a_n81_n597# a_n33_n500# w_n161_n600# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_5AQ4BN a_63_n500# a_n33_n500# a_n81_n597# w_n161_n620#
+ a_n125_n500#
X0 a_n33_n500# a_n81_n597# a_n125_n500# w_n161_n620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1 a_63_n500# a_n81_n597# a_n33_n500# w_n161_n620# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2 VPWR VGND A Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ZRN2GS a_n129_n500# a_63_n500# a_n225_n500# a_n321_n500#
+ a_n33_n500# a_n509_n500# a_n465_532# a_447_n500# a_159_n500# a_255_n500# a_351_n500#
+ a_n417_n500# VSUBS
X0 a_n417_n500# a_n465_532# a_n509_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X1 a_n33_n500# a_n465_532# a_n129_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X2 a_351_n500# a_n465_532# a_255_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X3 a_255_n500# a_n465_532# a_159_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X4 a_n321_n500# a_n465_532# a_n417_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X5 a_159_n500# a_n465_532# a_63_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X6 a_n225_n500# a_n465_532# a_n321_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X7 a_447_n500# a_n465_532# a_351_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X8 a_63_n500# a_n465_532# a_n33_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
X9 a_n129_n500# a_n465_532# a_n225_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_ZCCU26 a_n177_n1000# a_15_n1000# a_n269_n1000# a_207_n1000#
+ a_111_n1000# a_n81_n1000# a_n225_n1088# VSUBS
X0 a_207_n1000# a_n225_n1088# a_111_n1000# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X1 a_n177_n1000# a_n225_n1088# a_n269_n1000# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X2 a_111_n1000# a_n225_n1088# a_15_n1000# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X3 a_n81_n1000# a_n225_n1088# a_n177_n1000# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
X4 a_15_n1000# a_n225_n1088# a_n81_n1000# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+07u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_RPBXXN a_n33_n161# a_159_n161# a_n413_n161# a_255_n161#
+ w_n451_n269# a_n377_n258# a_351_n161# a_n129_n161# a_63_n161# a_n225_n161# a_n321_n161#
X0 a_255_n161# a_n377_n258# a_159_n161# w_n451_n269# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X1 a_n321_n161# a_n377_n258# a_n413_n161# w_n451_n269# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X2 a_159_n161# a_n377_n258# a_63_n161# w_n451_n269# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X3 a_n225_n161# a_n377_n258# a_n321_n161# w_n451_n269# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X4 a_63_n161# a_n377_n258# a_n33_n161# w_n451_n269# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X5 a_n129_n161# a_n377_n258# a_n225_n161# w_n451_n269# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X6 a_n33_n161# a_n377_n258# a_n129_n161# w_n451_n269# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
X7 a_351_n161# a_n377_n258# a_255_n161# w_n451_n269# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.61e+06u l=150000u
.ends

.subckt comparator VSS Vin_p Out_n Vin_n Out_p ext_clk VDD
Xx1 VSS VDD x2/A x1/A VSS VDD sky130_fd_sc_hd__buf_1
XXM13 x4/A x4/A x4/A x9/X VSS VSS VSS sky130_fd_pr__nfet_01v8_ZZU2YL
Xx2 VDD VSS x3/A x2/A VSS VDD sky130_fd_sc_hd__buf_4
Xx3 VSS VDD x3/A Out_p VSS VDD sky130_fd_sc_hd__buf_8
Xsky130_fd_pr__nfet_01v8_ZZU2YL_0 x1/A x1/A x1/A x4/A VSS VSS VSS sky130_fd_pr__nfet_01v8_ZZU2YL
Xx4 VSS VDD x5/A x4/A VSS VDD sky130_fd_sc_hd__buf_1
Xsky130_fd_pr__nfet_01v8_ZZU2YL_1 x4/A x4/A x4/A x1/A VSS VSS VSS sky130_fd_pr__nfet_01v8_ZZU2YL
Xx5 VDD VSS x6/A x5/A VSS VDD sky130_fd_sc_hd__buf_4
Xsky130_fd_pr__nfet_01v8_ZZU2YL_2 x1/A x1/A x1/A x9/X VSS VSS VSS sky130_fd_pr__nfet_01v8_ZZU2YL
Xx6 VSS VDD x6/A Out_n VSS VDD sky130_fd_sc_hd__buf_8
Xx7 VSS VDD x7/X ext_clk VSS VDD sky130_fd_sc_hd__buf_1
Xx8 VSS VDD x8/A x8/X VSS VDD sky130_fd_sc_hd__clkdlybuf4s15_1
Xx9 VDD VSS x9/X x9/A VSS VDD sky130_fd_sc_hd__buf_2
Xsky130_fd_pr__pfet_01v8_QPTUVJ_0 m1_11380_5940# m1_11380_5940# x1/A VDD m1_11380_5940#
+ VDD VDD sky130_fd_pr__pfet_01v8_QPTUVJ
XXM1 m1_12420_6100# VDD x16/X VDD m1_12420_6100# sky130_fd_pr__pfet_01v8_FBQ47L
Xsky130_fd_pr__pfet_01v8_QPTUVJ_1 m1_12240_5940# m1_12240_5940# x4/A VDD m1_12240_5940#
+ VDD VDD sky130_fd_pr__pfet_01v8_QPTUVJ
XXM2 m1_10470_6110# VDD x16/X VDD m1_10470_6110# sky130_fd_pr__pfet_01v8_5AQ4BN
Xsky130_fd_sc_hd__inv_2_0 VDD VSS x15/X x8/A VSS VDD sky130_fd_sc_hd__inv_2
XXM4 m1_10470_6110# m1_10470_6110# m1_9910_5690# m1_10470_6110# m1_9910_5690# m1_10470_6110#
+ Vin_n m1_10470_6110# m1_9910_5690# m1_10470_6110# m1_9910_5690# m1_9910_5690# VSS
+ sky130_fd_pr__nfet_01v8_ZRN2GS
XXM9 VSS VSS m1_9910_5690# VSS m1_9910_5690# m1_9910_5690# x15/X VSS sky130_fd_pr__nfet_01v8_ZCCU26
Xsky130_fd_pr__pfet_01v8_RPBXXN_0 x1/A x1/A x1/A m1_12240_5940# VDD m1_12420_6100#
+ x1/A m1_12240_5940# m1_12240_5940# x1/A m1_12240_5940# sky130_fd_pr__pfet_01v8_RPBXXN
Xsky130_fd_pr__nfet_01v8_ZRN2GS_0 m1_12420_6100# m1_12420_6100# m1_9910_5690# m1_12420_6100#
+ m1_9910_5690# m1_12420_6100# Vin_p m1_12420_6100# m1_9910_5690# m1_12420_6100# m1_9910_5690#
+ m1_9910_5690# VSS sky130_fd_pr__nfet_01v8_ZRN2GS
Xsky130_fd_pr__pfet_01v8_RPBXXN_1 x4/A x4/A x4/A m1_11380_5940# VDD m1_10470_6110#
+ x4/A m1_11380_5940# m1_11380_5940# x4/A m1_11380_5940# sky130_fd_pr__pfet_01v8_RPBXXN
Xx10 VSS VDD x8/X x11/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s15_1
Xx11 VSS VDD x11/A x9/A VSS VDD sky130_fd_sc_hd__clkdlybuf4s50_1
Xx12 VDD VSS x14/A x7/X VSS VDD sky130_fd_sc_hd__buf_2
Xx13 VDD VSS x15/X x16/A VSS VDD sky130_fd_sc_hd__inv_2
Xx14 VDD VSS x15/A x14/A VSS VDD sky130_fd_sc_hd__buf_4
Xx15 VSS VDD x15/A x15/X VSS VDD sky130_fd_sc_hd__buf_8
Xx16 VDD VSS x16/X x16/A VSS VDD sky130_fd_sc_hd__buf_4
.ends

.subckt all_analog V_in_p V_in_n comp_out_p sw_sample_unbuf comparator_clk sw_sp_n9
+ sw_sp_n8 sw_sp_n7 sw_sp_n6 sw_sp_n5 sw_sp_n4 sw_sp_n3 sw_sp_n2 sw_sp_n1 sw_sp_p9
+ sw_sp_p8 sw_sp_p7 sw_sp_p6 sw_sp_p5 sw_sp_p4 sw_sp_p3 sw_sp_p2 sw_sp_p1 sw_n8 sw_n7
+ sw_n6 sw_n5 sw_n4 sw_n3 sw_n2 sw_n1 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3 sw_p2 sw_p1
+ comp_out_n VDD VSS
Xdac_0 sw_sp_n9 sw_sp_n8 sw_sp_n7 sw_sp_n6 sw_sp_n5 sw_sp_n4 sw_sp_n3 sw_sp_n2 sw_sp_n1
+ sw_sp_p9 sw_sp_p8 sw_sp_p7 sw_sp_p6 sw_sp_p5 sw_sp_p4 sw_sp_p3 sw_sp_p2 sw_sp_p1
+ sw_n8 sw_n7 sw_n6 sw_n5 sw_n4 sw_n3 sw_n2 sw_n1 sw_p8 sw_p7 sw_p6 sw_p5 sw_p4 sw_p3
+ sw_p2 sw_p1 sw_sample_unbuf dac_0/sample_sw_buf_out VDD dac_0/Vin_p dac_0/Vin_n
+ VSS dac
Xsky130_fd_sc_hd__diode_2_0 VSS VDD sw_sp_p8 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_1 VSS VDD sw_sp_p6 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_2 VSS VDD sw_sp_p7 VDD VSS sky130_fd_sc_hd__diode_2
Xbootstrapped_sampling_switch_0 V_in_p V_in_n VDD VSS dac_0/sample_sw_buf_out dac_0/Vin_n
+ dac_0/Vin_p bootstrapped_sampling_switch
Xsky130_fd_sc_hd__diode_2_3 VSS VDD sw_sp_n6 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_4 VSS VDD sw_sp_n7 VDD VSS sky130_fd_sc_hd__diode_2
Xsky130_fd_sc_hd__diode_2_5 VSS VDD sw_sp_n8 VDD VSS sky130_fd_sc_hd__diode_2
Xcomparator_0 VSS dac_0/Vin_p comp_out_n dac_0/Vin_n comp_out_p comparator_clk VDD
+ comparator
.ends

.subckt sar_adc V_in_p V_in_n Done Clk Bit10 Bit9 Bit8 Bit7 Bit6 Bit5 Bit4 Bit3 Bit2
+ Bit1 RESET VDD VSS
Xcontroller_0 controller_0/sw_n1 controller_0/sw_n2 controller_0/sw_n3 controller_0/sw_n4
+ controller_0/sw_n5 controller_0/sw_n6 controller_0/sw_n7 controller_0/sw_n8 controller_0/sw_n_sp1
+ controller_0/sw_n_sp2 controller_0/sw_n_sp3 controller_0/sw_n_sp4 controller_0/sw_n_sp5
+ controller_0/sw_n_sp6 controller_0/sw_n_sp7 controller_0/sw_n_sp8 controller_0/sw_n_sp9
+ controller_0/sw_p1 controller_0/sw_p2 controller_0/sw_p3 controller_0/sw_p4 controller_0/sw_p5
+ controller_0/sw_p6 controller_0/sw_p7 controller_0/sw_p8 controller_0/sw_p_sp1 controller_0/sw_p_sp2
+ controller_0/sw_p_sp3 controller_0/sw_p_sp4 controller_0/sw_p_sp5 controller_0/sw_p_sp6
+ controller_0/sw_p_sp7 controller_0/sw_p_sp8 controller_0/sw_p_sp9 Bit1 Bit10 Bit2
+ Bit3 Bit4 Bit5 Bit6 Bit7 Bit8 Bit9 Clk controller_0/comp_out_n controller_0/comp_out_p
+ controller_0/comparator_clk Done RESET controller_0/sw_sample VDD VSS controller
Xall_analog_0 V_in_p V_in_n controller_0/comp_out_p controller_0/sw_sample controller_0/comparator_clk
+ controller_0/sw_n_sp9 controller_0/sw_n_sp8 controller_0/sw_n_sp7 controller_0/sw_n_sp6
+ controller_0/sw_n_sp5 controller_0/sw_n_sp4 controller_0/sw_n_sp3 controller_0/sw_n_sp2
+ controller_0/sw_n_sp1 controller_0/sw_p_sp9 controller_0/sw_p_sp8 controller_0/sw_p_sp7
+ controller_0/sw_p_sp6 controller_0/sw_p_sp5 controller_0/sw_p_sp4 controller_0/sw_p_sp3
+ controller_0/sw_p_sp2 controller_0/sw_p_sp1 controller_0/sw_n8 controller_0/sw_n7
+ controller_0/sw_n6 controller_0/sw_n5 controller_0/sw_n4 controller_0/sw_n3 controller_0/sw_n2
+ controller_0/sw_n1 controller_0/sw_p8 controller_0/sw_p7 controller_0/sw_p6 controller_0/sw_p5
+ controller_0/sw_p4 controller_0/sw_p3 controller_0/sw_p2 controller_0/sw_p1 controller_0/comp_out_n
+ VDD VSS all_analog
.ends

.subckt LNA_final Vgg_1v2 RF_in RF_out Vdd_1v8 Gnd
X0 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X3 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X5 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X11 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X12 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X13 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X15 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X16 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X21 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X24 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X25 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X26 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X27 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X28 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X29 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X31 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X33 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X34 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X37 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X38 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X41 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X42 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X45 a_n27544_n39610# a_n12387_n39359# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=1e+07u
X46 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X47 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X48 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X49 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X50 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X53 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X55 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X56 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X57 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X59 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X60 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X61 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X62 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X65 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X67 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X68 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X69 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X70 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
R0 Vgg_1v2 a_n27544_n39610# sky130_fd_pr__res_generic_po w=2e+06u l=1.053e+07u
X71 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X72 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X73 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X74 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X75 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X76 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X77 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X79 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X80 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X81 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X82 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X83 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X84 Gnd RF_out sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X85 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X86 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X87 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X88 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X89 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X90 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X91 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X92 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X93 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X94 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X95 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X96 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X97 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X98 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X99 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X100 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X102 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X103 Gnd RF_out sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X104 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X105 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X106 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X107 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X108 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X109 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X110 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X111 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X112 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X113 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X115 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X117 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X118 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X119 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X120 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X121 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X122 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X123 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X124 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X125 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X126 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X127 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X128 a_n12387_n39359# RF_in sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X129 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X130 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X131 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X132 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X133 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X134 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X135 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X136 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X137 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X138 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X139 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X140 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X141 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X142 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X143 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X144 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X145 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X146 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X147 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X148 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X149 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X150 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X151 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X152 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X153 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X154 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X155 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X156 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X157 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X158 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X159 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X160 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X161 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X162 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X163 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X164 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X165 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X166 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X167 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X168 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X169 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X170 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X171 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X172 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X173 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X174 Gnd Vdd_1v8 sky130_fd_pr__cap_mim_m3_2 l=1.5e+07u w=1.5e+07u
X175 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X176 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X177 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X178 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X179 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X180 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X181 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X182 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X183 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X184 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X185 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X186 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X187 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X188 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X189 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X190 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X191 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X192 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X193 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X194 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X195 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X196 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X197 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X198 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X199 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X200 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X201 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X202 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X203 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X204 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X205 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X206 a_38553_4766# Vdd_1v8 Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X207 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X208 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X209 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X210 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X211 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X212 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
D0 Gnd a_n12387_n39359# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X213 Vdd_1v8 Vdd_1v8 Vgg_1v2 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X214 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X215 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X216 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X217 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X218 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X219 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X220 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X221 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X222 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X223 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X224 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X225 Gnd Gnd Vgg_1v2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
D1 Gnd Vdd_1v8 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X226 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X227 Vgg_1v2 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X228 Vdd_1v8 Vdd_1v8 a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X229 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X230 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X231 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X232 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X233 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X234 Gnd Gnd Vdd_1v8 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X235 Gnd a_n12387_n39359# a_38553_4766# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X236 Vdd_1v8 Vdd_1v8 a_n27544_n39610# Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X237 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X238 Vgg_1v2 Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X239 a_n27544_n39610# Vdd_1v8 Vdd_1v8 Vdd_1v8 sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X240 a_38553_4766# a_n12387_n39359# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X241 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X242 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X243 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X244 Vdd_1v8 Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X245 a_n27544_n39610# Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X246 Gnd Gnd Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X247 Gnd Gnd a_n27544_n39610# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__res_high_po_2p85_DZGNGK a_3805_n2203# a_1351_n2203# a_5441_n2203#
+ a_n2739_n2203# a_n6829_n2203# a_n6829_1771# a_4623_1771# a_n4375_n2203# a_n4375_1771#
+ a_533_1771# a_n1103_n2203# a_6259_1771# a_2987_1771# a_n285_1771# a_n2739_1771#
+ a_5441_1771# a_2169_n2203# a_n6959_n2333# a_6259_n2203# a_4623_n2203# a_n5193_1771#
+ a_n1921_1771# a_n285_n2203# a_n3557_n2203# a_n1921_n2203# a_n5193_n2203# a_3805_1771#
+ a_2987_n2203# a_2169_1771# a_n3557_1771# a_1351_1771# a_n6011_n2203# a_533_n2203#
+ a_n1103_1771# a_n6011_1771#
X0 a_n5193_n2203# a_n5193_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X1 a_1351_n2203# a_1351_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X2 a_5441_n2203# a_5441_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X3 a_n2739_n2203# a_n2739_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X4 a_n6829_n2203# a_n6829_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X5 a_n1103_n2203# a_n1103_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X6 a_n3557_n2203# a_n3557_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X7 a_2169_n2203# a_2169_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X8 a_3805_n2203# a_3805_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X9 a_n285_n2203# a_n285_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X10 a_n6011_n2203# a_n6011_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X11 a_6259_n2203# a_6259_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X12 a_n1921_n2203# a_n1921_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X13 a_n4375_n2203# a_n4375_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X14 a_533_n2203# a_533_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X15 a_4623_n2203# a_4623_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X16 a_2987_n2203# a_2987_1771# a_n6959_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
.ends

.subckt r2r_8 vout b0 b1 b2 b3 b4 b5 b6 b7 vss
Xsky130_fd_pr__res_high_po_2p85_DZGNGK_0 b6 vss b7 b2 vss vss vss b1 m1_2567_4117#
+ m1_7475_4117# b3 vss vss vss m1_4203_4117# m1_12383_4117# b5 vss vss vss m1_931_8855#
+ vss vss m1_1749_143# vss m1_1749_143# m1_10747_4117# vss m1_9111_4117# vss vss b0
+ b4 m1_5839_4117# m1_931_4117# sky130_fd_pr__res_high_po_2p85_DZGNGK
Xsky130_fd_pr__res_high_po_2p85_DZGNGK_1 m1_10747_4117# m1_6657_8855# m1_12383_4117#
+ m1_4203_4117# vss vss vout m1_2567_4117# m1_1749_8855# m1_6657_8855# m1_5839_4117#
+ vss m1_9929_8855# m1_6657_8855# m1_3385_8855# vout m1_9111_4117# vss vss m1_9929_8855#
+ m1_1749_8855# m1_5021_8855# m1_5021_8855# m1_1749_8855# m1_3385_8855# m1_931_8855#
+ m1_9929_8855# m1_8293_8855# m1_8293_8855# m1_3385_8855# m1_8293_8855# m1_931_4117#
+ m1_7475_4117# m1_5021_8855# m1_931_8855# sky130_fd_pr__res_high_po_2p85_DZGNGK
.ends

.subckt sinv2_p a_n321_n70# a_n509_n70# w_n647_n289# a_n369_n167#
X0 a_n509_n70# a_n369_n167# a_n321_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n509_n70# a_n369_n167# a_n321_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n509_n70# a_n369_n167# a_n321_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n321_n70# a_n369_n167# a_n509_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n509_n70# a_n509_n70# a_n509_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n321_n70# a_n369_n167# a_n509_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X6 a_n509_n70# a_n509_n70# a_n509_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 a_n509_n70# a_n369_n167# a_n321_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X8 a_n321_n70# a_n369_n167# a_n509_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X9 a_n321_n70# a_n369_n167# a_n509_n70# w_n647_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt sinv2_n a_n419_n244# a_n177_92# a_n317_n70# a_n129_n70#
X0 a_n129_n70# a_n177_92# a_n317_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n317_n70# a_n177_92# a_n129_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n317_n70# a_n177_92# a_n129_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n317_n70# a_n317_n70# a_n317_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n317_n70# a_n317_n70# a_n317_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n129_n70# a_n177_92# a_n317_n70# a_n419_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt inv_simple2 m1_n42_n74# m2_584_n263# li_108_306# VSUBS
Xsinv2_p_0 m2_584_n263# li_108_306# li_108_306# m1_n42_n74# sinv2_p
Xsinv2_n_0 VSUBS m1_n42_n74# VSUBS m2_584_n263# sinv2_n
.ends

.subckt sinv_p w_n455_n289# a_n129_n70# a_n177_n167#
X0 w_n455_n289# a_n177_n167# a_n129_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 w_n455_n289# a_n177_n167# a_n129_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 w_n455_n289# w_n455_n289# w_n455_n289# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 w_n455_n289# w_n455_n289# w_n455_n289# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n129_n70# a_n177_n167# w_n455_n289# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n129_n70# a_n177_n167# w_n455_n289# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt sinv_n a_n81_92# a_n33_n70# a_n323_n244#
X0 a_n323_n244# a_n81_92# a_n33_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n33_n70# a_n81_92# a_n323_n244# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n323_n244# a_n323_n244# a_n323_n244# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n323_n244# a_n323_n244# a_n323_n244# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt inv_simple1 in out vdd vss
Xsinv_p_0 vdd out in sinv_p
Xsinv_n_0 in out vss sinv_n
.ends

.subckt inv_buffer2 in1 out1 vdd vss
Xinv_simple2_0 inv_simple1_0/out out1 vdd vss inv_simple2
Xinv_simple1_0 in1 inv_simple1_0/out vdd vss inv_simple1
.ends

.subckt slope_p a_n705_n70# a_591_n167# w_n1031_n289# a_15_n167# a_399_101# a_n753_101#
X0 w_n1031_n289# a_n753_101# a_n705_n70# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 w_n1031_n289# a_15_n167# a_n705_n70# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 w_n1031_n289# a_15_n167# a_n705_n70# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n705_n70# a_15_n167# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n705_n70# a_399_101# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 w_n1031_n289# a_399_101# a_n705_n70# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X6 w_n1031_n289# a_591_n167# a_n705_n70# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 w_n1031_n289# w_n1031_n289# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X8 a_n705_n70# a_591_n167# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X9 a_n705_n70# a_n753_101# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X10 w_n1031_n289# w_n1031_n289# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X11 a_n705_n70# a_n753_101# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X12 a_n705_n70# a_n753_101# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X13 w_n1031_n289# a_n753_101# a_n705_n70# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X14 w_n1031_n289# a_n753_101# a_n705_n70# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X15 a_n705_n70# a_n753_101# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X16 w_n1031_n289# a_n753_101# a_n705_n70# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X17 a_n705_n70# a_15_n167# w_n1031_n289# w_n1031_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt cap100f m3_n850_n800# c1_n750_n700#
X0 c1_n750_n700# m3_n850_n800# sky130_fd_pr__cap_mim_m3_1 l=7e+06u w=7e+06u
.ends

.subckt tg_p a_n221_n70# a_n33_n70# w_n359_n289# a_n81_101#
X0 a_n33_n70# a_n81_101# a_n221_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n221_n70# a_n221_n70# a_n221_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n221_n70# a_n221_n70# a_n221_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n221_n70# a_n81_101# a_n33_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt tg_n a_n221_n70# a_n33_n70# a_n323_n244# a_n81_n158#
X0 a_n221_n70# a_n81_n158# a_n33_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n33_n70# a_n81_n158# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n221_n70# a_n221_n70# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n221_n70# a_n221_n70# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt tg_1 sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289# sky130_fd_pr__pfet_01v8_X679XQ_0/a_n81_101#
+ sky130_fd_pr__nfet_01v8_2AA63J_0/a_n81_n158# m2_477_n333# m2_n53_n74# VSUBS
Xsky130_fd_pr__pfet_01v8_X679XQ_0 m2_477_n333# m2_n53_n74# sky130_fd_pr__pfet_01v8_X679XQ_0/w_n359_n289#
+ sky130_fd_pr__pfet_01v8_X679XQ_0/a_n81_101# tg_p
Xsky130_fd_pr__nfet_01v8_2AA63J_0 m2_477_n333# m2_n53_n74# VSUBS sky130_fd_pr__nfet_01v8_2AA63J_0/a_n81_n158#
+ tg_n
.ends

.subckt tgate_1 sw sw_out vdd vss sw_in
Xinv_simple1_0 sw inv_simple1_0/out vdd vss inv_simple1
Xtg_1_0 vdd sw inv_simple1_0/out sw_out sw_in vss tg_1
.ends

.subckt sinv_p2 a_n221_n70# a_n81_n167# a_n33_n70# w_n359_n289#
X0 a_n33_n70# a_n81_n167# a_n221_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n221_n70# a_n221_n70# a_n221_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n221_n70# a_n221_n70# a_n221_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n221_n70# a_n81_n167# a_n33_n70# w_n359_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt slopebuf bit1 bit0 bit2 clk_in clk_out vdd vbias vss
Xinv_buffer2_0 clk_in inv_simple1_0/in vdd vss inv_buffer2
Xinv_simple1_0 inv_simple1_0/in inv_simple1_0/out vdd vss inv_simple1
Xsky130_fd_pr__pfet_01v8_BDAFKN_0 m2_2652_919# vbias vdd tgate_1_2/sw_out tgate_1_1/sw_out
+ tgate_1_0/sw_out slope_p
Xcap100f_0 vss clk_out cap100f
Xsinv_n_0 inv_simple1_0/out clk_out vss sinv_n
Xtgate_1_1 bit0 tgate_1_1/sw_out vdd vss vbias tgate_1
Xtgate_1_0 bit2 tgate_1_0/sw_out vdd vss vbias tgate_1
Xtgate_1_2 bit1 tgate_1_2/sw_out vdd vss vbias tgate_1
Xsky130_fd_pr__pfet_01v8_X679XQ_0 m2_2652_919# inv_simple1_0/out clk_out vdd sinv_p2
.ends

.subckt sky130_fd_pr__res_high_po_2p85_97D7UQ a_7077_n2203# a_3805_n2203# a_1351_n2203#
+ a_5441_n2203# a_n2739_n2203# a_n6829_n2203# a_n6829_1771# a_4623_1771# a_n4375_n2203#
+ a_n8465_n2203# a_n4375_1771# a_533_1771# a_7895_n2203# a_7895_1771# a_n1103_n2203#
+ a_6259_1771# a_2987_1771# a_n285_1771# a_n2739_1771# a_n7647_1771# a_5441_1771#
+ a_2169_n2203# a_6259_n2203# a_4623_n2203# a_n8595_n2333# a_n5193_1771# a_n1921_1771#
+ a_n285_n2203# a_n3557_n2203# a_n1921_n2203# a_n5193_n2203# a_n7647_n2203# a_7077_1771#
+ a_3805_1771# a_2987_n2203# a_2169_1771# a_n3557_1771# a_n8465_1771# a_1351_1771#
+ a_n6011_n2203# a_533_n2203# a_n1103_1771# a_n6011_1771#
X0 a_n5193_n2203# a_n5193_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X1 a_1351_n2203# a_1351_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X2 a_5441_n2203# a_5441_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X3 a_n2739_n2203# a_n2739_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X4 a_n6829_n2203# a_n6829_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X5 a_7895_n2203# a_7895_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X6 a_n1103_n2203# a_n1103_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X7 a_n3557_n2203# a_n3557_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X8 a_n7647_n2203# a_n7647_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X9 a_2169_n2203# a_2169_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X10 a_3805_n2203# a_3805_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X11 a_n285_n2203# a_n285_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X12 a_n6011_n2203# a_n6011_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X13 a_6259_n2203# a_6259_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X14 a_n1921_n2203# a_n1921_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X15 a_n4375_n2203# a_n4375_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X16 a_n8465_n2203# a_n8465_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X17 a_533_n2203# a_533_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X18 a_4623_n2203# a_4623_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X19 a_7077_n2203# a_7077_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X20 a_2987_n2203# a_2987_1771# a_n8595_n2333# sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
.ends

.subckt r2r_10 b0 b1 b2 b3 b4 b5 b6 b7 vout b8 b9 vss
Xsky130_fd_pr__res_high_po_2p85_97D7UQ_0 m1_15655_4117# m1_12383_4117# m1_8293_8855#
+ m1_14019_4117# m1_5839_4117# m1_931_8855# m1_1749_8855# m1_13201_8855# m1_4203_4117#
+ vss m1_3385_8855# m1_8293_8855# vss vss m1_7475_4117# vout a_13201_4881# m1_8293_8855#
+ m1_5021_8855# m1_931_8855# m1_13201_8855# m1_10747_4117# m1_13201_8855# a_13201_4881#
+ vss m1_3385_8855# m1_6657_8855# m1_6657_8855# m1_3385_8855# m1_5021_8855# m1_1749_8855#
+ m1_931_4117# vout a_13201_4881# m1_9929_8855# m1_9929_8855# m1_5021_8855# vss m1_9929_8855#
+ m1_2567_4117# m1_9111_4117# m1_6657_8855# m1_1749_8855# sky130_fd_pr__res_high_po_2p85_97D7UQ
Xsky130_fd_pr__res_high_po_2p85_97D7UQ_1 b9 b7 vss b8 b3 m1_1749_143# m1_931_8855#
+ vss b2 vss m1_4203_4117# m1_9111_4117# vss vss b4 vss vss vss m1_5839_4117# m1_931_4117#
+ m1_14019_4117# b6 vss vss vss vss vss vss vss vss m1_1749_143# b0 m1_15655_4117#
+ m1_12383_4117# vss m1_10747_4117# vss vss vss b1 b5 m1_7475_4117# m1_2567_4117#
+ sky130_fd_pr__res_high_po_2p85_97D7UQ
.ends

.subckt sky130_fd_sc_hd__dfrtp_1$1 VGND VPWR Q RESET_B D CLK VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X13 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_2 VGND VPWR Q RESET_B D CLK VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X15 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X26 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt sky130_fd_sc_hd__decap_3$1 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_ef_sc_hd__decap_12$1 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt sky130_fd_sc_hd__decap_4$1 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__decap_6$1 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8$1 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__a221o_1 VPWR VGND X B1 A1 B2 A2 C1 VNB VPB
X0 a_465_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_109_297# B1 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_193_297# B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A2 a_193_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_193_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# B1 a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_297# C1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VGND A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_1$1 VGND VPWR X A VNB VPB
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=790000u l=150000u
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=520000u l=150000u
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR S A1 A0 X VNB VPB
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2_1 VGND VPWR A X B VNB VPB
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__conb_1$1 VGND VPWR LO HI VPB VNB
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_4$1 VGND VPWR X A VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__inv_2$1 VPWR VGND A Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3_1 VPWR VGND A X B C VNB VPB
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nor2_1 VGND VPWR B Y A VNB VPB
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_8 VGND VPWR X A VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or2b_1 VGND VPWR A B_N X VNB VPB
X0 a_219_297# a_27_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VGND B_N a_27_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR A a_301_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_219_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_301_297# a_27_53# a_219_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_219_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_27_53# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A a_219_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__buf_4$1 VPWR VGND X A VNB VPB
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xor2_1$1 VPWR VGND B X A VNB VPB
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2_1$1 VPWR VGND X B A VNB VPB
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__xnor2_1$1 VGND VPWR B Y A VNB VPB
X0 a_377_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_47_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_129_47# B a_47_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_285_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y a_47_47# a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A a_129_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_47_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_47_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Y B a_377_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1$1 VGND VPWR Y B A VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21oi_1 VPWR VGND A1 B1 Y A2 VNB VPB
X0 a_199_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_113_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR A1 a_113_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_113_297# B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A2 a_199_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a22o_1 VPWR VGND A1 A2 X B2 B1 VNB VPB
X0 VPWR A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_27_297# B1 a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A2 a_373_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_297# B1 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_373_47# A1 a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_109_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_109_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2111o_1 VGND VPWR B1 X D1 A1 A2 C1 VNB VPB
X0 VGND A2 a_660_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND C1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_414_297# C1 a_334_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND a_85_193# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_334_297# D1 a_85_193# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_516_297# B1 a_414_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_516_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_660_47# A1 a_85_193# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_85_193# D1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR A1 a_516_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_85_193# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR a_85_193# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2bb2a_1 VPWR VGND A1_N X A2_N B2 B1 VNB VPB
X0 a_206_369# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_206_369# A2_N a_205_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND B2 a_489_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_585_369# B2 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_47# a_206_369# a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_489_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR A2_N a_206_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_76_199# a_206_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_205_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR B1 a_585_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 VGND VPWR X A VNB VPB
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and2b_1 VGND VPWR X A_N B VNB VPB
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_1 VGND VPWR A2 A1 B1 Y VNB VPB
X0 Y A2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_27_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 a_109_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfstp_1$1 VPWR VGND D Q SET_B CLK VNB VPB
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X5 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X6 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=540000u l=150000u
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o221a_1 VGND VPWR A2 X B1 C1 A1 B2 VNB VPB
X0 a_240_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_51_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VGND A1 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_51_297# B2 a_245_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_149_47# C1 a_51_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_240_47# B1 a_149_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A1 a_512_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 X a_51_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_149_47# B2 a_240_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_245_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR C1 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_512_297# A2 a_51_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3b_1 VGND VPWR B C A_N Y VNB VPB
X0 Y a_53_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_232_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A_N a_53_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A_N a_53_93# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_316_47# B a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 Y a_53_93# a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o211a_1 VGND VPWR C1 B1 A2 A1 X VNB VPB
X0 VGND A1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_510_47# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_79_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_79_21# A2 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_297_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_79_21# C1 a_510_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_215_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and4_1 VGND VPWR X C A B D VNB VPB
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__and3_1 VGND VPWR X B A C VNB VPB
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 VPWR VGND Q CLK D VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a2bb2o_1 VGND VPWR B1 A1_N A2_N X B2 VNB VPB
X0 a_226_47# A2_N a_226_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_489_413# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_226_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR B2 a_489_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_489_413# a_226_47# a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_76_199# a_226_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VGND B1 a_556_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_556_47# B2 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VGND A2_N a_226_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 a_226_47# A1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__dfrtp_4$1 VGND VPWR Q RESET_B D CLK VNB VPB
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X12 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X16 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X17 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X18 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X29 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X30 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X31 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21boi_1 VPWR VGND Y A1 B1_N A2 VNB VPB
X0 a_300_297# a_27_413# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR A1 a_300_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_384_47# A1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 a_300_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1$1 VPWR VGND A X VNB VPB
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a32o_1 VGND VPWR X A3 B2 B1 A1 A2 VNB VPB
X0 a_93_21# A1 a_346_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_93_21# B1 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_584_47# B1 a_93_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_93_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND B2 a_584_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_256_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_250_297# B2 a_93_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND a_93_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_250_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A2 a_250_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_250_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_346_47# A2 a_256_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or3b_1 VGND VPWR A C_N X B VNB VPB
X0 a_109_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_215_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND a_109_93# a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VGND A a_215_53# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A a_369_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 a_369_297# B a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_215_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_297_297# a_109_93# a_215_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 X a_215_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o21ai_2 VGND VPWR B1 Y A2 A1 VNB VPB
X0 VGND A2 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 Y B1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_29_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y A2 a_112_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND A1 a_29_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_112_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_112_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_29_47# B1 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_29_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21o_1 VPWR VGND A2 A1 B1 X VNB VPB
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_4 VGND VPWR Y A B C VNB VPB
X0 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A a_445_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 a_27_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_445_47# A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X14 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_445_47# B a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VGND C a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a31o_1 VGND VPWR A2 B1 A1 A3 X VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__o31a_1 VGND VPWR X A2 B1 A1 A3 VNB VPB
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a41o_1 VGND VPWR A3 A4 A2 X B1 A1 VNB VPB
X0 a_465_47# A2 a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VGND A4 a_561_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A3 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_297_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_297_297# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A1 a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_381_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_297_297# B1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_79_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 a_561_47# A3 a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand3_1 VGND VPWR Y A C B VNB VPB
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_193_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y A a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_109_47# C VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22ai_1 VGND VPWR A2 B1 Y A1 B2 VNB VPB
X0 VGND A2 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_27_47# B2 Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 VPWR A1 a_307_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 a_307_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 a_27_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 Y B2 a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_109_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a211o_1 VGND VPWR X A2 B1 A1 C1 VNB VPB
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_80_21# C1 a_472_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A2 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_300_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 a_217_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_80_21# A1 a_300_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_472_297# B1 a_217_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_80_21# C1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o2111a_1 VPWR VGND X D1 C1 B1 A2 A1 VNB VPB
X0 a_676_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_512_47# B1 a_409_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_306_47# D1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VGND A2 a_512_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR C1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A1 a_676_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_512_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_409_47# C1 a_306_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_79_21# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__o22a_1 VGND VPWR A2 X B1 A1 B2 VNB VPB
X0 a_78_199# B1 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 VPWR A1 a_493_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 a_493_297# A2 a_78_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VPWR a_78_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A2 a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_78_199# B2 a_292_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_215_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 a_215_47# B2 a_78_199# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X8 a_292_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND a_78_199# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_fd_sc_hd__or4_1 VPWR VGND C A X B D VNB VPB
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__a21bo_1 VGND VPWR X A1 B1_N A2 VNB VPB
X0 a_298_297# a_27_413# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 a_215_297# a_27_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_298_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 VPWR B1_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_382_47# A1 a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 VGND B1_N a_27_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A1 a_298_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A2 a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt wrapper clk_in dac[0] dac[1] dac[2] dac[3] dac[4] dac[5] dac[6] dac[7] load
+ read ref_in reset s_in s_out vbias2[0] vbias2[1] vbias2[2] vbias2[3] vbias2[4] vbias2[5]
+ vbias2[6] vbias2[7] vco_in _0001_ _0002_ _0006_ _0010_ _0225_ _0226_ _0227_ _0229_
+ _0230_ _0463_ _0464_ _0470_ _0473_ _0480_ _0730_ _0732_ _0751_ _0752_ _0753_ _0754_
+ _0755_ _0757_ _0760_ _0798_ _0800_ _0912_ _0913_ _0914_ _0915_ _0918_ _0919_ _0920_
+ _0921_ _0923_ _0925_ _0930_ _0931_ _0932_ _0936_ _0938_ _0939_ _0940_ _0941_ _0942_
+ _0943_ d2.t_load\[13\] d2.t_load\[25\] d5.fll_core.counter1.count\[0\] d5.fll_core.counter1.count\[1\]
+ d5.fll_core.counter1.count\[2\] d5.fll_core.counter1.count\[4\] d5.fll_core.counter1.count\[5\]
+ d5.fll_core.counter1.count\[6\] d5.fll_core.counter1.count\[7\] d5.fll_core.counter1.count\[8\]
+ d5.fll_core.counter_reset net45 lock net6 net7 _0045_ _0146_ _0275_ _0276_ _0787_
+ _0788_ _0277_ _0278_ _0870_ _0875_ _0878_ _0881_ _0882_ _0883_ _0884_ _0885_ _0886_
+ _0888_ _0282_ _0381_ _0383_ _0384_ _0388_ _0389_ _0147_ _0148_ _0465_ _0467_ _0927_
+ _0468_ _0469_ _0149_ _0934_ _0150_ _0937_ _0151_ _0652_ _0671_ _0672_ _0673_ _0674_
+ clknet_4_15_0_clk_in d2.r_reg\[21\] d2.r_reg\[22\] d2.r_reg\[24\] d2.r_reg\[25\]
+ d2.r_reg\[27\] d2.r_reg\[28\] d2.r_reg\[31\] _0675_ d2.t_load\[19\] d2.t_load\[20\]
+ d2.t_load\[21\] d2.t_load\[23\] d2.t_load\[24\] _0677_ d2.t_load\[27\] d2.t_load\[28\]
+ d2.t_load\[30\] d2.t_load\[31\] _0678_ _0679_ _0681_ _0683_ _0684_ _0685_ _0686_
+ _0689_ _0154_ net44 _0158_ _0042_ _0043_ _0044_ _0700_ _0702_ _0704_ _0410_ _0412_
+ _0738_ _0739_ _0143_ _0267_ _0269_ _0271_ _0273_ clknet_4_12_0_clk_in clknet_4_13_0_clk_in
+ _0144_ d2.r_reg\[12\] d2.r_reg\[13\] d2.r_reg\[14\] d2.r_reg\[16\] d2.r_reg\[18\]
+ _0034_ _0773_ _0175_ _0176_ _0617_ _0177_ _0853_ d2.r_reg\[50\] d2.t_load\[10\]
+ d2.t_load\[11\] _0304_ d2.t_load\[15\] d2.t_load\[16\] d2.t_load\[17\] _0372_ _0373_
+ _0374_ _0375_ _0376_ _0377_ _0378_ _0379_ _0178_ _0889_ d2.t_load\[50\] d2.t_load\[51\]
+ _0890_ _0891_ _0894_ _0897_ _0040_ _0138_ _0139_ _0140_ _0690_ _0692_ _0694_ _0695_
+ _0696_ _0697_ _0698_ _0950_ _0952_ _0953_ _0956_ _0957_ _0958_ _0959_ _0960_ _0962_
+ _0965_ _0968_ clknet_0_ref_in clknet_1_1__leaf_ref_in _0509_ _0510_ _0513_ _0797_
+ _0514_ _0799_ _0515_ _0516_ _0518_ _0118_ _0120_ _0141_ _0457_ _0459_ _0462_ _0121_
+ _0124_ _0223_ _0000_ _0354_ _0355_ _0356_ d2.t_load\[18\] _0472_ _0358_ _0474_ _0475_
+ _0476_ _0477_ _0478_ _0359_ _0482_ _0485_ _0486_ _0487_ d5.fll_core.corner_tmp\[0\]
+ d5.fll_core.corner_tmp\[2\] _0488_ _0489_ _0490_ _0491_ _0492_ _0495_ _0496_ _0498_
+ _0502_ d5.fll_core.tmp\[0\] d5.fll_core.tmp\[1\] d5.fll_core.tmp\[3\] d5.fll_core.tmp\[6\]
+ _0504_ net43 _0506_ _0508_ _0945_ _0947_ _0948_ _0748_ _0749_ _0750_ _0777_ _0789_
+ _0859_ _0865_ _0866_ _0871_ _0872_ _0873_ _0874_ _0876_ _0877_ _0156_ _0880_ _0159_
+ _0286_ _0287_ _0288_ _0289_ _0290_ _0291_ _0640_ _0642_ clknet_4_11_0_clk_in _0644_
+ _0650_ _0651_ _0653_ _0654_ _0655_ _0657_ _0658_ _0661_ d2.r_reg\[29\] d2.r_reg\[30\]
+ _0662_ d2.r_reg\[32\] d2.r_reg\[33\] d2.r_reg\[34\] d2.r_reg\[36\] d2.r_reg\[37\]
+ d2.r_reg\[41\] _0663_ _0664_ _0665_ _0666_ _0669_ _0670_ vdd _0049_ _0050_ _0051_
+ d2.t_load\[29\] _0052_ d2.t_load\[33\] d2.t_load\[34\] d2.t_load\[39\] d2.t_load\[44\]
+ _0390_ _0391_ _0393_ _0394_ _0396_ _0400_ _0401_ _0402_ _0060_ net12 _0743_ _0164_
+ _0168_ _0630_ _0637_ _0864_ _0059_ _0641_ _0862_ d2.t_load\[36\] d2.t_load\[37\]
+ _0643_ d2.t_load\[41\] _0863_ _0868_ _0645_ d2.r_reg\[38\] _0646_ d2.r_reg\[42\]
+ _0647_ _0649_ _0292_ _0403_ _0293_ _0295_ _0297_ net17 net19 _0061_ _0163_ _0744_
+ net8 net9 _0745_ _0066_ _0593_ d2.t_load\[43\] d2.r_reg\[44\] _0595_ d2.r_reg\[61\]
+ d2.t_load\[62\] d2.r_reg\[62\] _0598_ _0629_ _0840_ _0635_ _0636_ _0083_ _0404_
+ _0405_ _0841_ _0296_ _0065_ _0187_ _0189_ _0424_ net26 net27 clknet_4_10_0_clk_in
+ _0315_ _0316_ _0317_ _0062_ clknet_4_8_0_clk_in _0302_ _0303_ _0071_ _0312_ _0313_
+ _0183_ _0184_ _0186_ _0855_ _0420_ _0190_ _0248_ _0249_ _0418_ _0171_ _0174_ _0172_
+ _0586_ _0790_ _0791_ _0250_ _0602_ d2.t_load\[45\] d2.t_load\[46\] _0604_ _0605_
+ d2.t_load\[57\] d2.t_load\[58\] d2.t_load\[60\] _0173_ _0618_ _0620_ _0622_ _0624_
+ _0626_ _0628_ _0079_ _0245_ _0631_ _0406_ _0409_ d5.fll_core.strobe d2.r_reg\[45\]
+ _0733_ _0734_ _0735_ d5.mux01.out\[3\] d5.mux01.out\[5\] d5.mux01.out\[6\] d5.mux01.out\[7\]
+ d2.r_reg\[46\] d2.r_reg\[47\] _0736_ d2.r_reg\[48\] d2.r_reg\[49\] _0633_ d2.r_reg\[51\]
+ d2.r_reg\[58\] _0737_ _0069_ _0417_ _0740_ _0070_ _0246_ _0247_ _0843_ _0300_ _0201_
+ _0202_ _0741_ _0742_ _0077_ _0588_ _0589_ _0308_ d2.r_reg\[54\] d2.r_reg\[55\] d2.r_reg\[56\]
+ _0310_ _0075_ d2.r_reg\[66\] d2.r_reg\[75\] _0836_ _0838_ _0414_ _0415_ _0076_ _0847_
+ _0849_ _0850_ _0851_ _0606_ _0607_ _0608_ _0609_ _0611_ _0086_ _0425_ d2.t_load\[54\]
+ d2.t_load\[55\] d2.t_load\[65\] _0435_ _0436_ _0320_ d5.fll_core.tmp\[9\] _0892_
+ d5.mux01.out\[9\] _0253_ _0181_ _0182_ _0095_ _0096_ _0192_ _0584_ _0585_ _0781_
+ _0782_ clknet_4_2_0_clk_in clknet_4_3_0_clk_in _0195_ _0590_ _0592_ _0792_ _0200_
+ _0594_ _0084_ _0085_ _0568_ _0569_ _0570_ _0571_ _0427_ _0429_ _0572_ _0434_ d2.r_reg\[63\]
+ _0579_ _0318_ _0319_ d2.r_reg\[68\] _0321_ _0323_ _0324_ d2.r_reg\[72\] _0581_ _0087_
+ _0825_ _0088_ _0089_ _0828_ _0094_ net23 net24 net25 _0833_ _0834_ _0582_ _0583_
+ _0839_ _0193_ _0194_ _0196_ _0433_ _0564_ _0091_ _0092_ _0197_ _0576_ net20 net21
+ net22 _0829_ _0830_ _0831_ _0832_ _0577_ _0578_ _0330_ d2.r_reg\[70\] _0431_ _0432_
+ _0559_ _0560_ _0561_ _0441_ _0442_ _0562_ clknet_4_1_0_clk_in _0203_ _0204_ _0563_
+ _0205_ _0566_ _0331_ _0332_ _0333_ _0793_ _0207_ _0334_ _0337_ _0104_ _0547_ _0548_
+ _0549_ _0550_ _0551_ _0817_ _0575_ _0552_ _0553_ _0554_ _0555_ _0556_ d2.r_reg\[77\]
+ d2.r_reg\[79\] d2.r_reg\[81\] net30 net31 net32 net33 _0819_ _0821_ _0098_ _0100_
+ _0101_ _0102_ _0824_ clknet_4_0_0_clk_in _0557_ _0453_ _0460_ _0973_ _0974_ _0976_
+ _0977_ _0980_ _0981_ _0984_ _0985_ _0986_ _0990_ _0991_ _0461_ _0761_ _0762_ _0763_
+ _0764_ _0765_ _0766_ _0768_ _0769_ _0785_ _0016_ _0011_ _0500_ _0501_ _0112_ _0528_
+ _0529_ _0532_ _0012_ _0013_ _0123_ _0015_ _0128_ _0236_ _0237_ _0240_ d5.fll_core.counter2.count\[1\]
+ d5.fll_core.counter2.count\[2\] d5.fll_core.counter2.count\[5\] d5.fll_core.counter2.count\[6\]
+ d5.fll_core.counter2.count\[7\] d5.fll_core.counter2.count\[8\] _0243_ _0244_ _0908_
+ net42 _0136_ _0137_ _0848_ _0264_ _0365_ d2.t_load\[3\] clknet_4_6_0_clk_in d2.t_load\[4\]
+ d2.t_load\[7\] d2.t_load\[8\] d2.t_load\[9\] _0306_ _0786_ _0366_ _0367_ _0368_
+ clknet_4_7_0_clk_in _0616_ _0025_ _0026_ _0030_ _0260_ _0073_ d2.r_reg\[4\] d2.r_reg\[5\]
+ d2.r_reg\[6\] d2.r_reg\[7\] d2.r_reg\[10\] _0129_ _0899_ _0901_ _0904_ d5.fll_core.tmp\[8\]
+ _0905_ _0259_ _0130_ d5.mux01.out\[8\] _0131_ _0179_ _0706_ _0708_ _0709_ _0710_
+ _0711_ _0712_ _0713_ _0714_ _0715_ _0716_ _0717_ _0718_ _0719_ _0720_ _0721_ _0722_
+ _0263_ _0134_ _0074_ d2.t_load\[1\] _0814_ _0530_ _0815_ _0774_ _0541_ _0542_ _0543_
+ _0544_ _0545_ _0546_ _0221_ _0816_ _0105_ net1 _0106_ _0349_ d2.r_reg\[84\] net2
+ d2.r_reg\[85\] _0256_ _0023_ _0802_ _0115_ _0783_ _0803_ _0211_ net28 _0212_ _0220_
+ _0519_ _0723_ net36 _0805_ _0725_ _0524_ _0806_ _0794_ _0255_ _0340_ _0116_ _0809_
+ _0810_ _0450_ _0811_ _0214_ _0216_ _0812_ _0813_ _0344_ _0521_ _0522_ _0362_ _0525_
+ _0526_ _0527_ _0909_ _0910_ _0795_ _0345_ _0347_ _0348_ _0108_ _0533_ _0534_ _0536_
+ net16 _0109_ _0537_ _0540_ _0451_ _0111_ _0350_ _0449_ d2.r_reg\[86\] d2.r_reg\[87\]
+ d2.r_reg\[88\] d2.r_reg\[89\] d2.r_reg\[90\] d2.t_load\[93\] d2.t_load\[94\] d2.r_reg\[93\]
+ d2.r_reg\[95\] d2.t_load\[0\] net39 net4 net40 _0456_ _0804_ _0728_ _0342_ _0127_
+ _0113_ _0114_ _0343_ _0447_ _0448_ corner[0] corner[1] corner[2] slope_ctrl[0] slope_ctrl[1]
+ slope_ctrl[2] vbias1[0] vbias1[1] vbias1[2] vbias1[3] vbias1[4] vbias1[5] vbias1[6]
+ vbias1[7] vbias3[0] vbias3[1] vbias3[2] vbias3[3] vbias3[4] vbias3[5] vbias3[6]
+ vbias3[7] _0003_ _0004_ _0005_ _0007_ _0008_ _0009_ _0228_ _0231_ _0232_ _0233_
+ _0234_ _0458_ _0731_ _0756_ _0758_ _0759_ _0911_ _0916_ _0917_ _0935_ clknet_0_vco_in
+ clknet_1_0__leaf_vco_in clknet_1_1__leaf_vco_in d5.fll_core.corner_tmp\[1\] d5.fll_core.counter1.count\[9\]
+ net5 _0682_ _0687_ _0688_ _0157_ _0041_ _0046_ _0047_ _0776_ _0879_ _0887_ _0152_
+ _0153_ _0279_ _0922_ _0924_ _0926_ _0928_ _0929_ _0933_ _0280_ clknet_0_clk_in _0281_
+ _0380_ _0382_ _0385_ _0386_ _0392_ d2.r_reg\[19\] d2.r_reg\[20\] d2.r_reg\[23\]
+ d2.r_reg\[26\] d2.t_load\[12\] d2.t_load\[22\] d2.t_load\[26\] _0155_ d5.fll_core.counter1.count\[3\]
+ _0466_ _0676_ _0680_ _0033_ _0142_ _0625_ _0268_ _0270_ _0272_ _0274_ _0145_ _0691_
+ _0693_ _0699_ _0701_ _0703_ _0705_ _0707_ _0035_ d2.r_reg\[11\] d2.r_reg\[15\] d2.r_reg\[17\]
+ _0036_ _0037_ _0038_ _0775_ d2.r_reg\[52\] _0039_ _0854_ _0031_ d2.t_load\[49\]
+ _0032_ _0895_ _0896_ _0898_ _0411_ _0483_ _0944_ _0946_ _0949_ _0951_ _0954_ _0955_
+ _0961_ _0963_ _0964_ _0966_ _0967_ _0969_ _0970_ _0971_ _0484_ _0493_ clknet_1_0__leaf_ref_in
+ _0494_ _0497_ _0499_ _0503_ _0505_ _0784_ _0796_ _0507_ _0511_ _0512_ _0517_ _0117_
+ _0119_ _0224_ d2.t_load\[14\] _0122_ _0125_ _0351_ _0352_ _0353_ _0471_ d5.fll_core.tmp\[2\]
+ d5.fll_core.tmp\[4\] d5.fll_core.tmp\[5\] d5.fll_core.tmp\[7\] _0479_ _0481_ _0747_
+ _0160_ _0161_ _0162_ _0387_ _0166_ _0395_ _0167_ _0048_ _0053_ _0054_ _0055_ _0056_
+ clknet_4_14_0_clk_in _0057_ _0627_ _0656_ _0659_ d2.r_reg\[35\] d2.r_reg\[39\] d2.r_reg\[40\]
+ _0660_ _0667_ _0668_ _0283_ d2.t_load\[32\] d2.t_load\[35\] d2.t_load\[40\] _0284_
+ d2.t_load\[56\] _0285_ _0294_ net13 net14 net15 _0638_ _0639_ _0648_ d2.t_load\[38\]
+ _0746_ d2.t_load\[42\] _0397_ _0867_ _0869_ _0398_ d2.r_reg\[43\] _0399_ net10 net11
+ _0165_ _0169_ _0058_ _0063_ _0423_ d2.t_load\[61\] _0596_ _0597_ _0298_ _0299_ _0599_
+ d2.r_reg\[60\] _0861_ _0170_ _0188_ _0634_ _0081_ _0082_ _0842_ _0778_ net18 _0421_
+ _0422_ _0064_ _0846_ _0600_ _0601_ _0603_ _0619_ _0621_ _0185_ d2.t_load\[47\] d2.t_load\[48\]
+ clknet_4_9_0_clk_in _0623_ d2.t_load\[59\] _0779_ d2.t_load\[63\] _0068_ _0632_
+ _0072_ _0078_ _0301_ _0305_ _0314_ d5.mux01.out\[0\] d5.mux01.out\[1\] d5.mux01.out\[2\]
+ d5.mux01.out\[4\] _0080_ _0856_ _0407_ _0251_ _0252_ _0408_ _0857_ _0419_ _0858_
+ d2.r_reg\[57\] d2.r_reg\[59\] _0860_ _0844_ _0845_ _0067_ _0826_ _0827_ _0835_ _0837_
+ _0311_ _0206_ _0416_ _0322_ _0610_ _0612_ _0613_ _0614_ _0325_ _0326_ d2.r_reg\[64\]
+ d2.r_reg\[65\] d2.r_reg\[67\] d2.r_reg\[69\] d2.r_reg\[71\] d2.r_reg\[73\] d2.r_reg\[74\]
+ d2.r_reg\[76\] d2.r_reg\[78\] d2.r_reg\[80\] d2.r_reg\[82\] d2.r_reg\[83\] _0327_
+ _0426_ _0428_ _0430_ _0437_ _0438_ _0439_ _0440_ _0443_ _0444_ _0328_ _0329_ _0335_
+ _0336_ _0338_ _0208_ d2.t_load\[64\] _0209_ _0210_ _0090_ _0093_ _0097_ _0180_ _0099_
+ _0103_ _0191_ _0198_ _0254_ _0558_ _0565_ _0567_ _0573_ _0574_ _0580_ _0587_ _0591_
+ _0780_ _0199_ _0309_ net29 net34 net35 _0818_ _0820_ _0822_ _0823_ _0360_ _0361_
+ _0363_ _0767_ _0770_ _0771_ _0531_ _0801_ _0807_ _0808_ _0019_ _0020_ d2.r_reg\[91\]
+ d2.r_reg\[92\] _0217_ _0218_ _0219_ _0903_ _0014_ _0017_ _0018_ d5.fll_core.counter2.count\[0\]
+ d5.fll_core.counter2.count\[3\] d5.fll_core.counter2.count\[4\] d5.fll_core.counter2.count\[9\]
+ _0235_ _0238_ _0452_ _0239_ _0241_ _0242_ _0126_ _0346_ _0972_ _0975_ net41 _0978_
+ _0979_ _0982_ _0983_ _0988_ _0989_ _0357_ _0906_ _0907_ _0029_ d2.t_load\[6\] _0265_
+ _0266_ _0135_ d2.r_reg\[3\] _0364_ _0024_ _0852_ _0027_ _0028_ d2.r_reg\[8\] _0369_
+ _0370_ d2.r_reg\[9\] _0413_ _0132_ d2.r_reg\[53\] _0133_ _0724_ _0726_ _0615_ d2.t_load\[2\]
+ _0371_ _0261_ _0893_ _0307_ _0900_ _0987_ d2.t_load\[52\] d2.t_load\[53\] _0902_
+ _0262_ _0258_ d2.t_load\[5\] _0446_ _0727_ net3 _0772_ _0454_ _0455_ d2.r_reg\[94\]
+ d2.r_reg\[2\] _0107_ clknet_4_4_0_clk_in d2.r_reg\[1\] _0339_ _0341_ _0729_ _0021_
+ _0022_ _0257_ _0445_ _0110_ d2.t_load\[95\] _0213_ _0535_ _0538_ _0523_ _0539_ _0222_
+ clknet_4_5_0_clk_in _0520_ net37 net38 _0215_ vss
X_2037_ vss vdd d2.r_reg\[32\] _0053_ _0287_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2106_ vss vdd d5.fll_core.tmp\[5\] _0122_ _0356_ clknet_1_1__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_39_277 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_52_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_22_111 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_22_177 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_45_269 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_45_247 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_45_203 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_26_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_36_258 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1270_ vdd vss _0982_ _0978_ d2.t_load\[1\] _0979_ _0977_ _0981_ vss vdd sky130_fd_sc_hd__a221o_1
X_1606_ vss vdd _0271_ _0695_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1537_ vss vdd _0630_ d2.t_load\[37\] d2.r_reg\[38\] _0648_ vss vdd sky130_fd_sc_hd__mux2_1
X_1468_ vss vdd _0596_ d2.r_reg\[59\] _0600_ _0601_ vss vdd sky130_fd_sc_hd__mux2_1
X_1399_ vss vdd _0336_ _0553_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_63_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_42_217 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_27_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_357 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_58_350 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_37_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_33_206 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_56_309 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1253_ vss vdd d5.fll_core.tmp\[5\] _0966_ d5.fll_core.tmp\[4\] vss vdd sky130_fd_sc_hd__or2_1
X_1322_ vss vdd _0491_ d5.fll_core.tmp\[7\] _0498_ _0499_ vss vdd sky130_fd_sc_hd__mux2_1
Xwrapper_44 vss vdd net44 wrapper_44/HI vdd vss sky130_fd_sc_hd__conb_1$1
XFILLER_64_353 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1184_ vss vdd _0904_ _0892_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_59_103 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_59_169 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_55_342 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_375 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_48_61 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_58_180 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_0_57 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_0_79 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1871_ vdd vss _0786_ _0139_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1940_ vdd vss _0793_ _0201_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_50_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1305_ vdd vss d5.fll_core.tmp\[9\] _0484_ d5.fll_core.tmp\[8\] d5.fll_core.tmp\[1\]
+ vss vdd sky130_fd_sc_hd__or3_1
X_1236_ vss vdd _0947_ _0949_ d5.fll_core.tmp\[8\] vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_52_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1098_ vss vdd _0407_ _0858_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1167_ vss vdd _0375_ _0895_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_37_386 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_12_209 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_60_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_264 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_161 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_43_356 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_43_345 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_34_96 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_34_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_50_62 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2070_ vss vdd d2.r_reg\[65\] _0086_ _0320_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1021_ vss vdd _0814_ d2.r_reg\[82\] net33 _0818_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_19_364 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1785_ vdd vss _0778_ _0061_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1923_ vdd vss _0791_ _0186_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1854_ vdd vss _0785_ _0123_ vss vdd sky130_fd_sc_hd__inv_2$1
Xclkbuf_4_6_0_clk_in vss vdd clknet_4_6_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
X_1219_ vss vdd d5.fll_core.counter1.count\[6\] d2.t_load\[26\] _0933_ vss vdd sky130_fd_sc_hd__or2b_1
X_2199_ vss vdd net39 _0215_ _0449_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_25_389 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_4_249 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_45_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_356 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_31_359 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1570_ vss vdd _0662_ d2.r_reg\[27\] _0670_ _0671_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_3_260 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_66_234 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2053_ vss vdd d2.r_reg\[48\] _0069_ _0303_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2122_ vss vdd d2.t_load\[11\] _0138_ _0372_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_34_197 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1004_ vss vdd _0803_ d2.r_reg\[90\] net41 _0809_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_19_194 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_22_326 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_22_348 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1768_ vdd vss _0776_ _0046_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1906_ vdd vss _0790_ _0780_ vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_30_370 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1837_ vdd vss _0783_ _0108_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1699_ vdd vss d5.fll_core.counter1.count\[0\] _0002_ d5.fll_core.counter1.count\[1\]
+ vss vdd sky130_fd_sc_hd__xor2_1$1
XFILLER_25_175 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_40_178 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_25_186 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_13_337 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_21_370 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xoutput7 vss vdd corner[2] net7 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput42 vss vdd vbias3[6] net42 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput20 vss vdd vbias1[0] net20 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput31 vss vdd vbias2[3] net31 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_0_230 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_48_278 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_63_248 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_131 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_153 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_16_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1622_ vss vdd _0706_ d2.r_reg\[11\] _0705_ _0707_ vss vdd sky130_fd_sc_hd__mux2_1
X_1553_ vss vdd _0652_ d2.t_load\[32\] d2.r_reg\[33\] _0659_ vss vdd sky130_fd_sc_hd__mux2_1
X_1484_ vss vdd _0596_ d2.r_reg\[54\] _0611_ _0612_ vss vdd sky130_fd_sc_hd__mux2_1
X_2036_ vss vdd d2.r_reg\[31\] _0052_ _0286_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2105_ vss vdd d5.fll_core.tmp\[4\] _0121_ _0355_ clknet_1_1__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_22_189 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_53_281 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_26_53 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_42_85 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_42_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_3_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_36_237 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_44_292 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1536_ vss vdd _0293_ _0647_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1605_ vss vdd _0684_ d2.r_reg\[16\] _0694_ _0695_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_59_318 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_59_307 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1467_ vss vdd _0586_ d2.t_load\[59\] d2.r_reg\[60\] _0600_ vss vdd sky130_fd_sc_hd__mux2_1
X_1398_ vss vdd _0552_ d2.r_reg\[81\] _0551_ _0553_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_42_229 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_2019_ vss vdd d2.r_reg\[14\] _0035_ _0269_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_18_237 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_53_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_26_292 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_174 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1252_ vdd vss _0965_ _0964_ _0963_ vss vdd sky130_fd_sc_hd__and2_1$1
X_1321_ vss vdd _0497_ _0498_ _0952_ vss vdd sky130_fd_sc_hd__xnor2_1$1
Xwrapper_45 vss vdd net45 wrapper_45/HI vdd vss sky130_fd_sc_hd__conb_1$1
XFILLER_64_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1183_ vss vdd _0367_ _0903_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_17_292 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_58_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1519_ vss vdd _0618_ d2.r_reg\[43\] _0635_ _0636_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_59_159 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_15_207 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_387 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_23_251 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_122 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_376 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_332 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1870_ vdd vss _0786_ _0138_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_9_89 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_43_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1304_ vss vdd _0483_ _0482_ _0947_ vss vdd sky130_fd_sc_hd__nand2_1$1
X_1166_ vss vdd _0893_ d2.r_reg\[14\] d2.t_load\[14\] _0895_ vss vdd sky130_fd_sc_hd__mux2_1
X_1235_ vdd vss _0948_ _0947_ d5.fll_core.tmp\[8\] vss vdd sky130_fd_sc_hd__and2_1$1
X_1097_ vss vdd _0848_ d2.r_reg\[46\] d2.t_load\[46\] _0858_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_20_221 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1999_ vdd vss _0795_ _0249_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_47_118 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_50_41 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_34_53 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_7_225 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1020_ vss vdd _0444_ _0817_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_19_321 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_198 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_187 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1922_ vdd vss _0791_ _0185_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_19_376 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1784_ vdd vss _0778_ _0773_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1853_ vdd vss _0785_ _0122_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_6_291 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1218_ vss vdd d5.fll_core.counter1.count\[5\] d2.t_load\[25\] _0932_ vss vdd sky130_fd_sc_hd__or2b_1
X_1149_ vss vdd _0383_ _0885_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_25_324 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2198_ vss vdd net38 _0214_ _0448_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_25_368 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_228 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_206 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_29_86 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_43_198 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_62 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_3_272 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2052_ vss vdd d2.r_reg\[47\] _0068_ _0302_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2121_ vss vdd d2.t_load\[10\] _0137_ _0371_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1003_ vss vdd _0452_ _0808_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1905_ vdd vss _0789_ _0170_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_30_382 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1767_ vdd vss _0776_ _0045_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1698_ vss vdd net15 _0750_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1836_ vdd vss _0783_ _0107_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_66_29 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_65_290 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_13_305 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_40_146 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_21_382 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
Xoutput10 vss vdd dac[2] net10 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput8 vss vdd dac[0] net8 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput43 vss vdd vbias3[7] net43 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput32 vss vdd vbias2[4] net32 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput21 vss vdd vbias1[1] net21 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_63_205 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_8_320 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_165 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1552_ vss vdd _0288_ _0658_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_8_353 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1621_ vss vdd _0706_ net1 vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_2104_ vss vdd d5.fll_core.tmp\[3\] _0120_ _0354_ clknet_1_1__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfrtp_2
X_1483_ vss vdd _0608_ d2.t_load\[54\] d2.r_reg\[55\] _0611_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_62_271 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2035_ vss vdd d2.r_reg\[30\] _0051_ _0285_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_22_124 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1819_ vdd vss _0782_ _0091_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_60_208 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_53_293 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_42_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_13_102 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_13_135 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_42_75 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_301 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_389 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_3_69 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_36_205 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_8_172 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1535_ vss vdd _0640_ d2.r_reg\[38\] _0646_ _0647_ vss vdd sky130_fd_sc_hd__mux2_1
X_1604_ vss vdd _0674_ d2.t_load\[16\] d2.r_reg\[17\] _0694_ vss vdd sky130_fd_sc_hd__mux2_1
X_1466_ vss vdd _0315_ _0599_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1397_ vss vdd _0552_ _0892_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_42_208 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2018_ vss vdd d2.r_reg\[13\] _0034_ _0268_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_35_271 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_12_56 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1320_ vdd vss _0951_ _0496_ _0497_ _0495_ vss vdd sky130_fd_sc_hd__a21oi_1
XFILLER_49_363 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1251_ vss vdd _0946_ _0964_ d5.fll_core.tmp\[4\] vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1182_ vss vdd _0893_ d2.r_reg\[6\] d2.t_load\[6\] _0903_ vss vdd sky130_fd_sc_hd__mux2_1
Xwrapper_46 vss vdd lock wrapper_46/HI vdd vss sky130_fd_sc_hd__conb_1$1
XFILLER_64_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_32_274 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_32_230 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_17_260 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_59_149 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1518_ vss vdd _0630_ d2.t_load\[43\] d2.r_reg\[44\] _0635_ vss vdd sky130_fd_sc_hd__mux2_1
X_1449_ vss vdd _0574_ d2.r_reg\[65\] _0587_ _0588_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_15_219 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_3_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_65_119 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_65_108 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_96 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_0_37 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_9_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1303_ vdd vss _0462_ d5.fll_core.counter1.count\[9\] _0482_ _0481_ _0480_ vss vdd
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_64_141 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_52_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1234_ vdd vss _0946_ _0947_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1096_ vss vdd _0408_ _0857_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1165_ vss vdd _0376_ _0894_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1998_ vdd vss _0795_ _0248_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_55_174 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_43_314 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_43_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_7_237 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_141 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_19_388 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1852_ vdd vss _0785_ _0121_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1921_ vdd vss _0791_ _0184_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_34_347 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1783_ vdd vss _0777_ _0060_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1217_ vss vdd _0928_ _0931_ _0930_ _0927_ d5.fll_core.counter1.count\[4\] _0929_
+ vss vdd sky130_fd_sc_hd__a2111o_1
X_1148_ vss vdd _0881_ d2.r_reg\[22\] d2.t_load\[22\] _0885_ vss vdd sky130_fd_sc_hd__mux2_1
X_1079_ vss vdd _0848_ d2.r_reg\[55\] _0847_ _0849_ vss vdd sky130_fd_sc_hd__mux2_1
X_2197_ vss vdd net37 _0213_ _0447_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_28_141 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_66_225 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2120_ vss vdd d2.t_load\[9\] _0136_ _0370_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_66_258 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2051_ vss vdd d2.r_reg\[46\] _0067_ _0301_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1002_ vss vdd _0803_ d2.r_reg\[91\] net42 _0808_ vss vdd sky130_fd_sc_hd__mux2_1
X_1904_ vdd vss _0789_ _0169_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1835_ vdd vss _0783_ _0106_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1766_ vdd vss _0776_ _0044_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1697_ vss vdd d2.t_load\[44\] d2.t_load\[41\] d2.t_load\[63\] _0750_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_57_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_136 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_114 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_21_350 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xoutput11 vss vdd dac[3] net11 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput9 vss vdd dac[1] net9 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_0_265 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xoutput33 vss vdd vbias2[5] net33 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput22 vss vdd vbias1[2] net22 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_56_280 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_56_85 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_56_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_31_125 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_177 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1551_ vss vdd _0640_ d2.r_reg\[33\] _0657_ _0658_ vss vdd sky130_fd_sc_hd__mux2_1
X_1620_ vss vdd _0696_ d2.t_load\[11\] d2.r_reg\[12\] _0705_ vss vdd sky130_fd_sc_hd__mux2_1
X_1482_ vss vdd _0310_ _0610_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_8_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2103_ vss vdd d5.fll_core.tmp\[2\] _0119_ _0353_ clknet_1_1__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_39_258 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_39_225 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_62_294 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2034_ vss vdd d2.r_reg\[29\] _0050_ _0284_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_22_136 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1818_ vdd vss _0782_ _0780_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1749_ vdd vss _0774_ _0029_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_26_66 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_42_65 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_13_169 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_42_98 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_357 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_3_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_66_3 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_8_184 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1534_ vss vdd _0630_ d2.t_load\[38\] d2.r_reg\[39\] _0646_ vss vdd sky130_fd_sc_hd__mux2_1
X_1603_ vss vdd _0272_ _0693_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1465_ vss vdd _0596_ d2.r_reg\[60\] _0598_ _0599_ vss vdd sky130_fd_sc_hd__mux2_1
X_2017_ vss vdd d2.r_reg\[12\] _0033_ _0267_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1396_ vss vdd _0542_ net32 d2.r_reg\[82\] _0551_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_50_253 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_10_106 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_2_305 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_26_261 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_286 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_121 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_165 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_49_342 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1250_ vss vdd _0946_ _0963_ d5.fll_core.tmp\[5\] vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1181_ vss vdd _0368_ _0902_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_24_209 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_64_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1517_ vss vdd _0299_ _0634_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1448_ vss vdd _0586_ d2.t_load\[65\] d2.r_reg\[66\] _0587_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_55_356 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1379_ vss vdd _0342_ _0539_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_2_157 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_2_135 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_53 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_46_345 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_323 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_0_49 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_64_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_61_359 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_61_326 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_14_275 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1302_ vdd vss _0477_ _0481_ d2.t_load\[18\] d5.fll_core.counter1.count\[9\] _0462_
+ vss vdd sky130_fd_sc_hd__o2bb2a_1
X_1233_ vss vdd _0946_ _0945_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_29_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_64_197 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1095_ vss vdd _0848_ d2.r_reg\[47\] d2.t_load\[47\] _0857_ vss vdd sky130_fd_sc_hd__mux2_1
X_1164_ vss vdd _0893_ d2.r_reg\[15\] d2.t_load\[15\] _0894_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_37_323 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1997_ vdd vss _0795_ _0247_ vss vdd sky130_fd_sc_hd__inv_2$1
Xclkbuf_4_11_0_clk_in vss vdd clknet_4_11_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
Xclkbuf_0_clk_in vss vdd clknet_0_clk_in clk_in vss vdd sky130_fd_sc_hd__clkbuf_16
XFILLER_28_378 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_7_249 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_34_337 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1920_ vdd vss _0791_ _0183_ vss vdd sky130_fd_sc_hd__inv_2$1
Xclkbuf_1_0__f_ref_in vss vdd clknet_1_0__leaf_ref_in clknet_0_ref_in vss vdd sky130_fd_sc_hd__clkbuf_16
X_1851_ vdd vss _0785_ _0780_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1782_ vdd vss _0777_ _0059_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1216_ vss vdd _0930_ d2.t_load\[25\] d5.fll_core.counter1.count\[5\] vss vdd sky130_fd_sc_hd__and2b_1
XFILLER_37_142 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2196_ vss vdd net36 _0212_ _0446_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1147_ vss vdd _0384_ _0884_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1078_ vss vdd _0848_ _0802_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_25_359 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_25_337 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_25_315 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_25_304 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_1_81 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_45_65 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_43_123 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_28_197 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_28_131 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_66_248 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2050_ vss vdd d2.r_reg\[45\] _0066_ _0300_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_10_90 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_34_156 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1001_ vss vdd _0453_ _0807_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1765_ vdd vss _0776_ _0043_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1903_ vdd vss _0789_ _0168_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_30_340 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1834_ vdd vss _0783_ _0105_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1696_ vss vdd net14 _0749_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_65_281 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_25_101 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2179_ vss vdd net19 _0195_ _0429_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_15_68 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xoutput12 vss vdd dac[4] net12 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput34 vss vdd vbias2[6] net34 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput23 vss vdd vbias1[3] net23 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_0_277 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_56_292 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_56_53 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_16_189 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_8_333 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_8_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_12_351 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1550_ vss vdd _0652_ d2.t_load\[33\] d2.r_reg\[34\] _0657_ vss vdd sky130_fd_sc_hd__mux2_1
X_1481_ vss vdd _0596_ d2.r_reg\[55\] _0609_ _0610_ vss vdd sky130_fd_sc_hd__mux2_1
X_2033_ vss vdd d2.r_reg\[28\] _0049_ _0283_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_47_281 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2102_ vss vdd d5.fll_core.tmp\[1\] _0118_ _0352_ clknet_1_1__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_11_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1748_ vdd vss _0774_ _0028_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1817_ vdd vss _0781_ _0090_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1679_ vss vdd _0847_ d2.t_load\[53\] d5.fll_core.tmp\[8\] _0741_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_38_292 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_13_148 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_21_181 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_3_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_5_314 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_369 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_36_229 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_59_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1602_ vss vdd _0684_ d2.r_reg\[17\] _0692_ _0693_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_8_141 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1533_ vss vdd _0294_ _0645_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1464_ vss vdd _0586_ d2.t_load\[60\] d2.r_reg\[61\] _0598_ vss vdd sky130_fd_sc_hd__mux2_1
X_1395_ vss vdd _0337_ _0550_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2016_ vss vdd d2.r_reg\[11\] _0032_ _0266_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_50_298 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_10_118 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_12_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_58_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_58_343 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_221 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_1_361 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_64_346 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1180_ vss vdd _0893_ d2.r_reg\[7\] d2.t_load\[7\] _0902_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_17_273 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_32_298 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1516_ vss vdd _0618_ d2.r_reg\[44\] _0633_ _0634_ vss vdd sky130_fd_sc_hd__mux2_1
Xclkbuf_4_9_0_clk_in vss vdd clknet_4_9_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
X_1447_ vss vdd _0586_ _0519_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1378_ vss vdd _0530_ d2.r_reg\[87\] _0538_ _0539_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_23_57 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_64_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_58_173 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_357 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_9_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_14_221 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_14_298 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1301_ vss vdd _0476_ _0472_ _0479_ _0480_ vss vdd sky130_fd_sc_hd__o21ai_1
X_1232_ vss vdd _0945_ _0944_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_49_195 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1094_ vss vdd _0409_ _0856_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_37_379 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1163_ vss vdd _0893_ _0892_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1996_ vdd vss _0795_ _0246_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_55_187 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_36_390 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_11_257 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_50_55 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_59_97 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_61_146 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_124 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1781_ vdd vss _0777_ _0058_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1850_ vdd vss _0784_ _0120_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_41_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1215_ vss vdd _0929_ d2.t_load\[26\] d5.fll_core.counter1.count\[6\] vss vdd sky130_fd_sc_hd__and2b_1
X_1146_ vss vdd _0881_ d2.r_reg\[23\] d2.t_load\[23\] _0884_ vss vdd sky130_fd_sc_hd__mux2_1
X_2195_ vss vdd net35 _0211_ _0445_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_52_157 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_33_371 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1077_ vss vdd _0847_ d2.t_load\[55\] vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_1_93 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1979_ vdd vss _0800_ _0230_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_20_69 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_45_88 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_43_135 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_43_113 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_16_305 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_51_190 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_20_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_19_165 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1000_ vss vdd _0803_ d2.r_reg\[92\] net43 _0807_ vss vdd sky130_fd_sc_hd__mux2_1
X_1902_ vdd vss _0789_ _0167_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_34_146 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_22_319 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1764_ vdd vss _0776_ _0042_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1833_ vdd vss _0783_ _0104_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1695_ vss vdd d2.t_load\[44\] d2.t_load\[40\] d2.t_load\[62\] _0749_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_65_271 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1129_ vss vdd _0870_ d2.r_reg\[31\] d2.t_load\[31\] _0875_ vss vdd sky130_fd_sc_hd__mux2_1
X_2178_ vss vdd net18 _0194_ _0428_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_2
XFILLER_25_124 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
Xoutput13 vss vdd dac[5] net13 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_31_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xoutput24 vss vdd vbias1[4] net24 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput35 vss vdd vbias2[7] net35 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_48_249 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_0_245 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XPHY_130 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_31_138 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_24_190 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_8_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1480_ vss vdd _0608_ d2.t_load\[55\] d2.r_reg\[56\] _0609_ vss vdd sky130_fd_sc_hd__mux2_1
X_2032_ vss vdd d2.r_reg\[27\] _0048_ _0282_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2101_ vdd vss _0351_ d5.fll_core.tmp\[0\] _0117_ clknet_1_1__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfstp_1$1
XFILLER_30_182 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1678_ vss vdd d5.mux01.out\[7\] _0740_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1816_ vdd vss _0781_ _0089_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1747_ vdd vss _0774_ _0027_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_7_81 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_53_252 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_53_241 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_45_219 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_26_79 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_109 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_21_193 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_3_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_5_348 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_44_285 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1532_ vss vdd _0640_ d2.r_reg\[39\] _0644_ _0645_ vss vdd sky130_fd_sc_hd__mux2_1
X_1601_ vss vdd _0674_ d2.t_load\[17\] d2.r_reg\[18\] _0692_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_8_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1463_ vss vdd _0316_ _0597_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1394_ vss vdd _0530_ d2.r_reg\[82\] _0549_ _0550_ vss vdd sky130_fd_sc_hd__mux2_1
X_2015_ vss vdd d2.r_reg\[10\] _0031_ _0265_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_12_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_58_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_41_200 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_26_285 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_189 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_5_134 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_1_373 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1515_ vss vdd _0630_ d2.t_load\[44\] d2.r_reg\[45\] _0633_ vss vdd sky130_fd_sc_hd__mux2_1
X_1446_ vss vdd _0321_ _0585_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1377_ vss vdd _0520_ net38 d2.r_reg\[88\] _0538_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_23_299 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_23_69 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_64_65 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_61_317 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_58_152 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_0_29 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1300_ vss vdd _0477_ _0479_ _0473_ _0478_ d2.t_load\[18\] d2.t_load\[17\] vss vdd
+ sky130_fd_sc_hd__o221a_1
X_1231_ vdd vss _0944_ _0943_ _0940_ vss vdd sky130_fd_sc_hd__and2_1$1
XFILLER_37_347 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_37_303 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1162_ vss vdd _0892_ net1 vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_64_155 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_52_317 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1093_ vss vdd _0848_ d2.r_reg\[48\] d2.t_load\[48\] _0856_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_45_380 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1995_ vdd vss _0795_ _0245_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1429_ vdd vss _0574_ _0892_ vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_28_358 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_28_347 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_58 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_11_203 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_11_225 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_46_122 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_169 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_42_372 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_42_361 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1780_ vdd vss _0777_ _0057_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_34_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1145_ vss vdd _0385_ _0883_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1214_ vss vdd _0928_ d2.t_load\[27\] d5.fll_core.counter1.count\[7\] vss vdd sky130_fd_sc_hd__and2b_1
XFILLER_52_125 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_37_199 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_37_155 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2194_ vss vdd net34 _0210_ _0444_ clknet_4_1_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1076_ vss vdd _0417_ _0846_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1978_ vdd vss _0800_ _0229_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_29_79 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_29_68 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_29_57 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_51_180 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_10_70 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_13_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1901_ vdd vss _0789_ _0166_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1832_ vdd vss _0783_ _0103_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1694_ vss vdd net13 _0748_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1763_ vdd vss _0776_ _0041_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1128_ vss vdd _0393_ _0874_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1059_ vss vdd _0836_ d2.r_reg\[64\] d2.t_load\[64\] _0838_ vss vdd sky130_fd_sc_hd__mux2_1
X_2177_ vss vdd net17 _0193_ _0427_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_25_169 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_15_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xoutput14 vss vdd dac[6] net14 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput25 vss vdd vbias1[5] net25 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_31_69 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
Xoutput36 vss vdd vbias3[0] net36 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_0_202 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_206 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_131 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_120 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_8_346 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2100_ vss vdd d2.r_reg\[95\] _0116_ _0350_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_62_264 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2031_ vss vdd d2.r_reg\[26\] _0047_ _0281_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_54_209 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_0 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1815_ vdd vss _0781_ _0088_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1677_ vss vdd _0847_ d2.t_load\[52\] d5.fll_core.tmp\[7\] _0740_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_7_93 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1746_ vdd vss _0774_ _0026_ vss vdd sky130_fd_sc_hd__inv_2$1
X_2229_ vss vdd d5.fll_core.counter2.count\[7\] _0242_ _0018_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_5_327 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1531_ vss vdd _0630_ d2.t_load\[39\] d2.r_reg\[40\] _0644_ vss vdd sky130_fd_sc_hd__mux2_1
X_1600_ vss vdd _0273_ _0691_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1462_ vss vdd _0596_ d2.r_reg\[61\] _0595_ _0597_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_32_90 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_8_165 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1393_ vss vdd _0542_ net33 d2.r_reg\[83\] _0549_ vss vdd sky130_fd_sc_hd__mux2_1
X_2014_ vss vdd d2.r_reg\[9\] _0030_ _0264_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1729_ vss vdd _0767_ _0016_ _0766_ vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_58_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_37_57 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_26_231 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_18_209 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_53_67 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_113 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_64_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1514_ vss vdd _0300_ _0632_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1445_ vss vdd _0574_ d2.r_reg\[66\] _0584_ _0585_ vss vdd sky130_fd_sc_hd__mux2_1
X_1376_ vss vdd _0343_ _0537_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_23_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_48_67 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_307 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_58_197 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_9_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1230_ vss vdd _0936_ _0942_ _0916_ _0943_ vss vdd sky130_fd_sc_hd__nand3b_1
XFILLER_49_142 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1161_ vss vdd _0377_ _0891_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1092_ vss vdd _0410_ _0855_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1994_ vdd vss _0801_ _0244_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_9_293 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_28_304 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1428_ vss vdd _0564_ net22 d2.r_reg\[72\] _0573_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_18_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_43_329 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1359_ vss vdd _0904_ d2.r_reg\[93\] _0525_ _0526_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_11_237 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_11_215 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_59_77 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_46_156 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_19_304 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_19_337 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_61_159 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_137 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1213_ vdd vss d2.t_load\[24\] _0927_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1144_ vss vdd _0881_ d2.r_reg\[24\] d2.t_load\[24\] _0883_ vss vdd sky130_fd_sc_hd__mux2_1
X_1075_ vss vdd _0836_ d2.r_reg\[56\] d2.t_load\[56\] _0846_ vss vdd sky130_fd_sc_hd__mux2_1
X_2193_ vss vdd net33 _0209_ _0443_ clknet_4_1_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_18_370 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1977_ vdd vss _0800_ _0228_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_45_57 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_43_159 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_28_167 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_6_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_281 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_34_115 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_19_145 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1900_ vdd vss _0789_ _0165_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1831_ vdd vss _0783_ _0102_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_15_362 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1693_ vss vdd d2.t_load\[44\] d2.t_load\[39\] d2.t_load\[61\] _0748_ vss vdd sky130_fd_sc_hd__mux2_1
X_1762_ vdd vss _0776_ _0773_ vss vdd sky130_fd_sc_hd__buf_4$1
X_2176_ vss vdd d2.t_load\[65\] _0192_ _0426_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1127_ vss vdd _0870_ d2.r_reg\[32\] d2.t_load\[32\] _0874_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_40_129 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_107 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_33_181 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1058_ vss vdd _0426_ _0837_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_15_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_31_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xoutput15 vss vdd dac[7] net15 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput26 vss vdd vbias1[6] net26 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_0_258 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xoutput37 vss vdd vbias3[1] net37 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_56_273 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_132 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_121 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_110 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_31_118 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_12_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2030_ vss vdd d2.r_reg\[25\] _0046_ _0280_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XPHY_1 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1814_ vdd vss _0781_ _0087_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1745_ vdd vss _0774_ _0025_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1676_ vss vdd d5.mux01.out\[6\] _0739_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2159_ vss vdd d2.t_load\[48\] _0175_ _0409_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2228_ vss vdd d5.fll_core.counter2.count\[6\] _0241_ _0017_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_53_276 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_265 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1530_ vss vdd _0295_ _0643_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1461_ vss vdd _0596_ _0892_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1392_ vss vdd _0338_ _0548_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2013_ vss vdd d2.r_reg\[8\] _0029_ _0263_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_50_279 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_50_235 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_35_254 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1728_ vdd vss d5.fll_core.counter2.count\[4\] d5.fll_core.counter2.count\[5\] _0767_
+ _0763_ vss vdd sky130_fd_sc_hd__a21oi_1
XFILLER_2_309 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1659_ vss vdd d2.t_load\[33\] d2.t_load\[31\] d5.fll_core.corner_tmp\[1\] _0731_
+ vss vdd sky130_fd_sc_hd__mux2_1
Xclkbuf_4_14_0_clk_in vss vdd clknet_4_14_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
XFILLER_53_57 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_5_103 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_158 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_32_202 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_57_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1513_ vss vdd _0618_ d2.r_reg\[45\] _0631_ _0632_ vss vdd sky130_fd_sc_hd__mux2_1
X_1444_ vss vdd _0564_ net17 d2.r_reg\[67\] _0584_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_4_180 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1375_ vss vdd _0530_ d2.r_reg\[88\] _0536_ _0537_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_63_371 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_349 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_316 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_23_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_58_187 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_58_121 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_22_290 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_1_194 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_64_179 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_64_135 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1160_ vss vdd _0881_ d2.r_reg\[16\] d2.t_load\[16\] _0891_ vss vdd sky130_fd_sc_hd__mux2_1
X_1091_ vss vdd _0848_ d2.r_reg\[49\] d2.t_load\[49\] _0855_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_37_316 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1993_ vdd vss _0801_ _0243_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_9_261 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_227 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_124 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1358_ vss vdd _0520_ d2.t_load\[93\] d2.r_reg\[94\] _0525_ vss vdd sky130_fd_sc_hd__mux2_1
X_1427_ vss vdd _0327_ _0572_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1289_ vss vdd d2.t_load\[10\] _0001_ _0467_ d2.t_load\[11\] _0468_ vss vdd sky130_fd_sc_hd__o211a_1
XFILLER_36_382 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_34_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_50_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_11_249 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_59_89 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_46_135 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_6_253 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1212_ vss vdd _0926_ _0924_ _0922_ _0923_ _0925_ vss vdd sky130_fd_sc_hd__and4_1
X_2192_ vss vdd net32 _0208_ _0442_ clknet_4_0_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1143_ vss vdd _0386_ _0882_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1074_ vss vdd _0418_ _0845_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_37_135 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_360 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_382 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1976_ vdd vss _0800_ _0227_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_29_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_28_157 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xclkbuf_4_2_0_clk_in vss vdd clknet_4_2_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
XFILLER_66_208 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_19_124 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_19_157 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1761_ vdd vss _0775_ _0040_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1830_ vdd vss _0783_ _0101_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_15_374 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1692_ vss vdd net12 _0747_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1126_ vss vdd _0394_ _0873_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2175_ vss vdd d2.t_load\[64\] _0191_ _0425_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_33_193 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1057_ vss vdd _0836_ d2.r_reg\[65\] d2.t_load\[65\] _0837_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_15_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_21_333 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_31_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1959_ vdd vss _0794_ _0219_ vss vdd sky130_fd_sc_hd__inv_2$1
Xoutput27 vss vdd vbias1[7] net27 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput16 vss vdd s_out net16 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_0_215 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xoutput38 vss vdd vbias3[2] net38 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XPHY_100 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_133 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_122 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_111 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_31_108 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_12_300 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_12_322 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_12_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_230 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_62_211 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_296 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_2 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1813_ vdd vss _0781_ _0086_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_7_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_7_370 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1744_ vdd vss _0774_ _0024_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1675_ vss vdd _0847_ d2.t_load\[51\] d5.fll_core.tmp\[6\] _0739_ vss vdd sky130_fd_sc_hd__mux2_1
X_1109_ vss vdd _0402_ _0864_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_53_200 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2158_ vss vdd d2.t_load\[47\] _0174_ _0408_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2227_ vss vdd d5.fll_core.counter2.count\[5\] _0240_ _0016_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2089_ vss vdd d2.r_reg\[84\] _0105_ _0339_ clknet_4_1_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_42_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_44_233 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_29_274 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_16_60 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_12_163 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1460_ vss vdd _0586_ d2.t_load\[61\] d2.r_reg\[62\] _0595_ vss vdd sky130_fd_sc_hd__mux2_1
X_1391_ vss vdd _0530_ d2.r_reg\[83\] _0547_ _0548_ vss vdd sky130_fd_sc_hd__mux2_1
X_2012_ vss vdd d2.r_reg\[7\] _0028_ _0262_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1658_ vss vdd net5 _0730_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1727_ vss vdd _0766_ d5.fll_core.counter2.count\[5\] d5.fll_core.counter2.count\[4\]
+ _0763_ vss vdd sky130_fd_sc_hd__and3_1
XFILLER_12_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_58_314 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1589_ vss vdd _0684_ _0892_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_37_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_41_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_32_258 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_27_92 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_17_299 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1512_ vss vdd _0630_ d2.t_load\[45\] d2.r_reg\[46\] _0631_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_55_306 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1443_ vss vdd _0322_ _0583_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_4_170 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_85 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_4_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1374_ vss vdd _0520_ net39 d2.r_reg\[89\] _0536_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_63_383 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_23_236 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_23_225 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_23_258 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_23_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_58_166 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1090_ vss vdd _0411_ _0854_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_54_90 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1992_ vdd vss _0801_ _0242_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_9_273 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_55_136 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_103 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1288_ vdd vss d5.fll_core.counter1.count\[1\] _0467_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1357_ vss vdd _0349_ _0524_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1426_ vss vdd _0552_ d2.r_reg\[72\] _0571_ _0572_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_36_372 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_50_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_46_147 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_34_309 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_42_386 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_6_221 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_6_265 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1211_ vss vdd d5.fll_core.counter1.count\[8\] d2.t_load\[28\] _0925_ vss vdd sky130_fd_sc_hd__or2b_1
X_1142_ vss vdd _0881_ d2.r_reg\[25\] d2.t_load\[25\] _0882_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_1_20 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2191_ vss vdd net31 _0207_ _0441_ clknet_4_0_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_52_106 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1073_ vss vdd _0836_ d2.r_reg\[57\] d2.t_load\[57\] _0845_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_33_364 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_33_342 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_33_331 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1975_ vdd vss _0800_ _0226_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_20_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_29_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1409_ vss vdd _0542_ net28 d2.r_reg\[78\] _0560_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_45_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_16_309 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_61_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_150 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_34_128 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_27_180 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_15_342 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_15_386 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_19_169 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1691_ vss vdd d2.t_load\[44\] d2.t_load\[38\] d2.t_load\[60\] _0747_ vss vdd sky130_fd_sc_hd__mux2_1
X_1760_ vdd vss _0775_ _0039_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_32_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1125_ vss vdd _0870_ d2.r_reg\[33\] d2.t_load\[33\] _0873_ vss vdd sky130_fd_sc_hd__mux2_1
X_2174_ vss vdd d2.t_load\[63\] _0190_ _0424_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_33_161 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1056_ vss vdd _0836_ _0802_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_21_312 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1889_ vdd vss _0788_ _0155_ vss vdd sky130_fd_sc_hd__inv_2$1
Xoutput17 vss vdd slope_ctrl[0] net17 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_31_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xoutput28 vss vdd vbias2[0] net28 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput39 vss vdd vbias3[3] net39 vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1958_ vdd vss _0794_ _0218_ vss vdd sky130_fd_sc_hd__inv_2$1
XPHY_123 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_56_264 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XPHY_112 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_101 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_12_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_62_278 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_30_131 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_120 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XPHY_3 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_15_183 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1674_ vss vdd d5.mux01.out\[5\] _0738_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1812_ vdd vss _0781_ _0085_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_7_382 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1743_ vdd vss _0774_ _0023_ vss vdd sky130_fd_sc_hd__inv_2$1
X_2226_ vss vdd d5.fll_core.counter2.count\[4\] _0239_ _0015_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1108_ vss vdd _0859_ d2.r_reg\[41\] d2.t_load\[41\] _0864_ vss vdd sky130_fd_sc_hd__mux2_1
X_2157_ vss vdd d2.t_load\[46\] _0173_ _0407_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_38_253 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1039_ vss vdd _0435_ _0827_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2088_ vss vdd d2.r_reg\[83\] _0104_ _0338_ clknet_4_1_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_44_278 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_94 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_12_175 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_12_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1390_ vss vdd _0542_ net34 d2.r_reg\[84\] _0547_ vss vdd sky130_fd_sc_hd__mux2_1
X_2011_ vss vdd d2.r_reg\[6\] _0027_ _0261_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_50_248 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1657_ vss vdd d2.t_load\[33\] d2.t_load\[30\] d5.fll_core.corner_tmp\[0\] _0730_
+ vss vdd sky130_fd_sc_hd__mux2_1
X_1588_ vss vdd _0674_ d2.t_load\[21\] d2.r_reg\[22\] _0683_ vss vdd sky130_fd_sc_hd__mux2_1
X_1726_ vss vdd _0763_ _0015_ _0765_ vss vdd sky130_fd_sc_hd__xnor2_1$1
X_2209_ vdd vss d5.fll_core.corner_tmp\[0\] clknet_1_1__leaf_ref_in _0457_ vss vdd
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_53_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_64_318 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_40_270 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1511_ vss vdd _0630_ net2 vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1442_ vss vdd _0574_ d2.r_reg\[67\] _0582_ _0583_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_4_193 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_48_370 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_97 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_4_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1373_ vss vdd _0344_ _0535_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1709_ vss vdd _0756_ _0006_ _0755_ vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_48_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_58_134 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_13_73 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_60_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_60_354 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_62_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_13_292 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1991_ vdd vss _0801_ _0241_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1425_ vss vdd _0564_ net23 d2.r_reg\[73\] _0571_ vss vdd sky130_fd_sc_hd__mux2_1
X_1287_ vdd vss d5.fll_core.counter1.count\[2\] _0466_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_28_318 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1356_ vss vdd _0904_ d2.r_reg\[94\] _0523_ _0524_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_18_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_63_181 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_50_49 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_59_69 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_42_354 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_42_343 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_6_233 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_40_93 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1210_ vss vdd d5.fll_core.counter1.count\[9\] d2.t_load\[29\] _0924_ vss vdd sky130_fd_sc_hd__or2b_1
X_1141_ vss vdd _0881_ _0802_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1072_ vss vdd _0419_ _0844_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2190_ vss vdd net30 _0206_ _0440_ clknet_4_1_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_1_32 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_18_340 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1974_ vdd vss _0800_ _0225_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_29_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1408_ vss vdd _0333_ _0559_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1339_ vss vdd _0491_ d5.fll_core.tmp\[3\] _0511_ _0512_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_45_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_36_181 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_24_365 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_3_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_10_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_262 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1690_ vss vdd net11 _0746_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_25_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1124_ vss vdd _0395_ _0872_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2173_ vss vdd d2.t_load\[62\] _0189_ _0423_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1055_ vss vdd _0427_ _0835_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_18_170 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1957_ vdd vss _0794_ _0217_ vss vdd sky130_fd_sc_hd__inv_2$1
Xoutput18 vss vdd slope_ctrl[1] net18 vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1888_ vdd vss _0788_ _0154_ vss vdd sky130_fd_sc_hd__inv_2$1
Xoutput29 vss vdd vbias2[1] net29 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_56_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XPHY_124 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_113 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_102 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_16_118 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_21_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_21_73 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_47_243 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1811_ vdd vss _0781_ _0084_ vss vdd sky130_fd_sc_hd__inv_2$1
XPHY_4 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_15_195 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1673_ vss vdd _0847_ d2.t_load\[50\] d5.fll_core.tmp\[5\] _0738_ vss vdd sky130_fd_sc_hd__mux2_1
X_1742_ vdd vss _0774_ _0022_ vss vdd sky130_fd_sc_hd__inv_2$1
X_2225_ vss vdd d5.fll_core.counter2.count\[3\] _0238_ _0014_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1107_ vss vdd _0403_ _0863_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2156_ vss vdd d2.t_load\[45\] _0172_ _0406_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2087_ vss vdd d2.r_reg\[82\] _0103_ _0337_ clknet_4_1_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1038_ vss vdd _0825_ d2.r_reg\[74\] net25 _0827_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_29_254 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_8_136 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_12_187 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_4_331 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2010_ vss vdd d2.r_reg\[5\] _0026_ _0260_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_50_205 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1725_ vdd vss d5.fll_core.counter2.count\[4\] _0765_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_58_305 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1587_ vss vdd _0277_ _0682_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1656_ vss vdd _0255_ _0729_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2139_ vss vdd d2.t_load\[28\] _0155_ _0389_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2208_ vdd vss _0000_ d5.fll_core.counter_reset _0224_ clknet_1_1__leaf_ref_in vss
+ vdd sky130_fd_sc_hd__dfstp_1$1
XFILLER_37_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_53_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_34_290 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_49_305 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_32_238 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_43_82 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1510_ vss vdd _0301_ _0629_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1441_ vss vdd _0564_ net18 d2.r_reg\[68\] _0582_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_4_65 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1372_ vss vdd _0530_ d2.r_reg\[89\] _0534_ _0535_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_23_205 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1708_ vdd vss d5.fll_core.counter1.count\[4\] d5.fll_core.counter1.count\[5\] _0756_
+ _0753_ vss vdd sky130_fd_sc_hd__a21oi_1
X_1639_ vss vdd _0519_ d2.t_load\[5\] d2.r_reg\[6\] _0718_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_66_190 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_64_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_1_142 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_60_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_60_300 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1990_ vdd vss _0801_ _0240_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_13_260 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_9_286 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1355_ vss vdd _0520_ d2.t_load\[94\] d2.r_reg\[95\] _0523_ vss vdd sky130_fd_sc_hd__mux2_1
X_1424_ vss vdd _0328_ _0570_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1286_ vdd vss d5.fll_core.counter1.count\[3\] _0465_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_36_341 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_36_330 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xclkbuf_1_1__f_vco_in vss vdd clknet_1_1__leaf_vco_in clknet_0_vco_in vss vdd sky130_fd_sc_hd__clkbuf_16
XFILLER_51_333 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_34_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_1_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_6_245 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1140_ vss vdd _0387_ _0880_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1071_ vss vdd _0836_ d2.r_reg\[58\] d2.t_load\[58\] _0844_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_1_44 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_60_163 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1973_ vdd vss _0800_ d5.fll_core.counter_reset vss vdd sky130_fd_sc_hd__buf_4$1
X_1338_ vss vdd _0510_ _0511_ _0954_ vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1407_ vss vdd _0552_ d2.r_reg\[78\] _0558_ _0559_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_45_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_43_108 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_171 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1269_ vss vdd _0980_ d2.t_load\[1\] _0977_ _0981_ d2.t_load\[7\] vss vdd sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_10_53 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_34_108 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_19_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_19_138 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_42_163 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_347 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_15_333 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_15_355 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_71 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_65_211 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2172_ vss vdd d2.t_load\[61\] _0188_ _0422_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2241_ vss vdd d2.t_load\[65\] _0254_ d5.mux01.out\[9\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
XFILLER_2_270 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_18_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1123_ vss vdd _0870_ d2.r_reg\[34\] d2.t_load\[34\] _0872_ vss vdd sky130_fd_sc_hd__mux2_1
X_1054_ vss vdd _0825_ d2.r_reg\[66\] net17 _0835_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_18_182 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1887_ vdd vss _0788_ _0153_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_33_174 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1956_ vdd vss _0794_ _0216_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_21_358 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xoutput19 vss vdd slope_ctrl[2] net19 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XPHY_125 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_114 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_103 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_24_130 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_47_211 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_62_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_5 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_15_141 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1810_ vdd vss _0781_ _0083_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_11_380 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1741_ vdd vss _0774_ _0021_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1672_ vss vdd d5.mux01.out\[4\] _0737_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1106_ vss vdd _0859_ d2.r_reg\[42\] d2.t_load\[42\] _0863_ vss vdd sky130_fd_sc_hd__mux2_1
X_2155_ vss vdd d2.t_load\[44\] _0171_ _0405_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_4$1
XFILLER_38_277 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2224_ vss vdd d5.fll_core.counter2.count\[2\] _0237_ _0013_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_53_225 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_42_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2086_ vss vdd d2.r_reg\[81\] _0102_ _0336_ clknet_4_0_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1037_ vss vdd _0436_ _0826_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1939_ vdd vss _0793_ _0772_ vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_44_258 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_12_100 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_74 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_16_85 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_4_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_35_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_35_236 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1724_ vss vdd _0764_ _0014_ _0763_ vss vdd sky130_fd_sc_hd__nor2_1
X_1586_ vss vdd _0662_ d2.r_reg\[22\] _0681_ _0682_ vss vdd sky130_fd_sc_hd__mux2_1
X_1655_ vss vdd _0802_ net16 _0728_ _0729_ vss vdd sky130_fd_sc_hd__mux2_1
X_2138_ vss vdd d2.t_load\[27\] _0154_ _0388_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2207_ vss vdd d5.fll_core.strobe _0223_ _0000_ clknet_1_1__leaf_ref_in vss vdd sky130_fd_sc_hd__dfrtp_4$1
X_2069_ vss vdd d2.r_reg\[64\] _0085_ _0319_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_53_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_57_361 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_49_317 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_17_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_283 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_4_77 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1371_ vss vdd _0520_ net40 d2.r_reg\[90\] _0534_ vss vdd sky130_fd_sc_hd__mux2_1
X_1440_ vss vdd _0323_ _0581_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_23_217 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1707_ vss vdd _0755_ d5.fll_core.counter1.count\[4\] d5.fll_core.counter1.count\[5\]
+ _0753_ vss vdd sky130_fd_sc_hd__and3_1
X_1638_ vss vdd _0261_ _0717_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1569_ vss vdd _0652_ d2.t_load\[27\] d2.r_reg\[28\] _0670_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_46_309 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
Xclkbuf_4_5_0_clk_in vss vdd clknet_4_5_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
XFILLER_13_20 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_49_169 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_45_353 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_20_209 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1285_ vdd vss d5.fll_core.counter1.count\[4\] _0464_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_48_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1354_ vss vdd _0350_ _0522_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1423_ vss vdd _0552_ d2.r_reg\[73\] _0569_ _0570_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_51_345 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_48_180 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_367 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_50_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_42_334 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_24_52 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_24_41 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_24_96 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_10_253 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_10_286 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_27_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_60_131 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1070_ vss vdd _0420_ _0843_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_18_353 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1972_ vss vdd _0459_ _0799_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_33_378 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1337_ vdd vss _0510_ d5.fll_core.tmp\[2\] _0509_ _0947_ vss vdd sky130_fd_sc_hd__a21boi_1
X_1268_ vdd vss d5.fll_core.counter2.count\[7\] _0980_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1406_ vss vdd _0542_ net29 d2.r_reg\[79\] _0558_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_61_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1199_ vss vdd _0912_ _0913_ _0911_ vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_35_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_19_96 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_359 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_326 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_30_315 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1122_ vss vdd _0396_ _0871_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2171_ vss vdd d2.t_load\[60\] _0187_ _0421_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2240_ vss vdd d2.t_load\[64\] _0253_ d5.mux01.out\[8\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
XFILLER_2_282 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1053_ vss vdd _0428_ _0834_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_21_326 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_21_337 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1886_ vdd vss _0788_ _0152_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1955_ vdd vss _0794_ _0215_ vss vdd sky130_fd_sc_hd__inv_2$1
XPHY_126 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_115 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_104 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_24_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_12_359 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_47_256 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_6 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_15_153 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1671_ vss vdd _0847_ d2.t_load\[49\] d5.fll_core.tmp\[4\] _0737_ vss vdd sky130_fd_sc_hd__mux2_1
X_1740_ vdd vss _0774_ _0773_ vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_7_330 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_7_363 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_53_215 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1105_ vss vdd _0404_ _0862_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2154_ vss vdd d2.t_load\[43\] _0170_ _0404_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2223_ vss vdd d5.fll_core.counter2.count\[1\] _0236_ _0012_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2085_ vss vdd d2.r_reg\[80\] _0101_ _0335_ clknet_4_0_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_61_281 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1036_ vss vdd _0825_ d2.r_reg\[75\] net26 _0826_ vss vdd sky130_fd_sc_hd__mux2_1
X_1869_ vdd vss _0786_ _0137_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1938_ vdd vss _0792_ _0200_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_29_289 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_29_267 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_53 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_32_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_4_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_57_93 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1723_ vss vdd _0761_ _0764_ d5.fll_core.counter2.count\[3\] vss vdd sky130_fd_sc_hd__nor2_1
X_1654_ vss vdd _0519_ d2.t_load\[0\] d2.r_reg\[1\] _0728_ vss vdd sky130_fd_sc_hd__mux2_1
X_1585_ vss vdd _0674_ d2.t_load\[22\] d2.r_reg\[23\] _0681_ vss vdd sky130_fd_sc_hd__mux2_1
X_2206_ vss vdd d2.t_load\[95\] _0222_ _0456_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2137_ vss vdd d2.t_load\[26\] _0153_ _0387_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2068_ vss vdd d2.r_reg\[63\] _0084_ _0318_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1019_ vss vdd _0814_ d2.r_reg\[83\] net34 _0817_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_57_373 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_43_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_240 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_295 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_4_152 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1370_ vss vdd _0345_ _0533_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1706_ vss vdd _0753_ _0005_ _0464_ vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1637_ vss vdd _0706_ d2.r_reg\[6\] _0716_ _0717_ vss vdd sky130_fd_sc_hd__mux2_1
X_1568_ vss vdd _0283_ _0669_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_48_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1499_ vss vdd _0608_ d2.t_load\[49\] d2.r_reg\[50\] _0622_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_54_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_13_32 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_8_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_64_107 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_45_387 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_13_240 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1422_ vss vdd _0564_ net24 d2.r_reg\[74\] _0569_ vss vdd sky130_fd_sc_hd__mux2_1
X_1284_ vdd vss d5.fll_core.counter1.count\[5\] _0463_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1353_ vss vdd _0904_ d2.r_reg\[95\] _0521_ _0522_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_51_379 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_51_313 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_0999_ vss vdd _0454_ _0806_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_59_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_27_387 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_27_310 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_42_379 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_10_221 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_40_85 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_40_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_37_107 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_65_93 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_33_357 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_33_324 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_1_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_18_321 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_60_187 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1971_ vss vdd _0796_ d5.fll_core.corner_tmp\[2\] _0946_ _0799_ vss vdd sky130_fd_sc_hd__mux2_1
X_1405_ vss vdd _0334_ _0557_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1198_ vss vdd _0912_ d2.t_load\[23\] d5.fll_core.counter1.count\[3\] vss vdd sky130_fd_sc_hd__and2b_1
X_1336_ vss vdd _0509_ _0960_ _0955_ vss vdd sky130_fd_sc_hd__nand2_1$1
X_1267_ vss vdd d2.t_load\[9\] _0979_ d5.fll_core.counter2.count\[9\] vss vdd sky130_fd_sc_hd__or2_1
XFILLER_28_107 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xinput1 vdd vss load net1 vss vdd sky130_fd_sc_hd__dlymetal6s2s_1$1
XFILLER_59_276 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_10_77 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_15_313 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_84 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xclkbuf_0_vco_in vss vdd clknet_0_vco_in vco_in vss vdd sky130_fd_sc_hd__clkbuf_16
X_1121_ vss vdd _0870_ d2.r_reg\[35\] d2.t_load\[35\] _0871_ vss vdd sky130_fd_sc_hd__mux2_1
X_2170_ vss vdd d2.t_load\[59\] _0186_ _0420_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1052_ vss vdd _0825_ d2.r_reg\[67\] net18 _0834_ vss vdd sky130_fd_sc_hd__mux2_1
X_1954_ vdd vss _0794_ _0214_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_21_305 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1885_ vdd vss _0788_ _0151_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_56_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XPHY_116 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_105 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1319_ vdd vss _0496_ _0947_ d5.fll_core.tmp\[6\] vss vdd sky130_fd_sc_hd__and2_1$1
XPHY_127 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_12_338 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_21_98 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_95 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_146 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_7 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_15_165 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1670_ vss vdd d5.mux01.out\[3\] _0736_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2222_ vss vdd d5.fll_core.counter2.count\[0\] _0235_ _0011_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_23_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2153_ vss vdd d2.t_load\[42\] _0169_ _0403_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1104_ vss vdd _0859_ d2.r_reg\[43\] d2.t_load\[43\] _0862_ vss vdd sky130_fd_sc_hd__mux2_1
X_1035_ vss vdd _0825_ _0802_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_2084_ vss vdd d2.r_reg\[79\] _0100_ _0334_ clknet_4_0_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1937_ vdd vss _0792_ _0199_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_21_113 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_21_146 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1868_ vdd vss _0786_ _0136_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1799_ vdd vss _0779_ _0074_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_52_293 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_52_271 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_249 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_32_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_4_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_345 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1584_ vss vdd _0278_ _0680_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1722_ vdd vss _0763_ _0761_ d5.fll_core.counter2.count\[3\] vss vdd sky130_fd_sc_hd__and2_1$1
X_1653_ vss vdd _0256_ _0727_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_66_330 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2205_ vss vdd d2.t_load\[94\] _0221_ _0455_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2136_ vss vdd d2.t_load\[25\] _0152_ _0386_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_41_208 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2067_ vss vdd d2.r_reg\[62\] _0083_ _0317_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1018_ vss vdd _0445_ _0816_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_1_337 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_57_385 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_57_330 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_27_20 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_17_205 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_25_260 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_197 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_0_370 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_16_282 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1705_ vss vdd _0754_ _0004_ _0753_ vss vdd sky130_fd_sc_hd__nor2_1
X_1567_ vss vdd _0662_ d2.r_reg\[28\] _0668_ _0669_ vss vdd sky130_fd_sc_hd__mux2_1
X_1636_ vss vdd _0696_ d2.t_load\[6\] d2.r_reg\[7\] _0716_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_64_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1498_ vss vdd _0305_ _0621_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2119_ vss vdd d2.t_load\[8\] _0135_ _0369_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_54_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_13_44 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_38_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_60_347 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_54_62 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_38_96 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_13_274 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1421_ vss vdd _0329_ _0568_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1283_ vdd vss d2.t_load\[19\] _0462_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1352_ vss vdd _0520_ d2.t_load\[95\] net4 _0521_ vss vdd sky130_fd_sc_hd__mux2_1
X_0998_ vss vdd _0803_ d2.r_reg\[93\] d2.t_load\[93\] _0806_ vss vdd sky130_fd_sc_hd__mux2_1
X_1619_ vss vdd _0267_ _0704_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_54_152 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_42_325 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_20 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_24_76 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_10_233 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_10_266 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_40_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_49_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_1_69 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1970_ vss vdd _0458_ _0798_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_45_152 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_53_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1335_ vss vdd _0355_ _0508_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_5_281 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1404_ vss vdd _0552_ d2.r_reg\[79\] _0556_ _0557_ vss vdd sky130_fd_sc_hd__mux2_1
X_1197_ vss vdd _0911_ d2.t_load\[22\] d5.fll_core.counter1.count\[2\] vss vdd sky130_fd_sc_hd__and2b_1
XFILLER_36_163 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1266_ vss vdd _0978_ d5.fll_core.counter2.count\[9\] d2.t_load\[9\] vss vdd sky130_fd_sc_hd__nand2_1$1
XFILLER_24_314 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xinput2 vss vdd net2 read vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_3_218 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_42_188 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_2_295 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_65_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1120_ vss vdd _0870_ _0802_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1051_ vss vdd _0429_ _0833_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1884_ vdd vss _0788_ _0780_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1953_ vdd vss _0794_ _0213_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_56_236 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1318_ vdd vss _0947_ _0966_ _0495_ _0965_ _0962_ vss vdd sky130_fd_sc_hd__a22o_1
XPHY_128 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_117 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_106 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1249_ vss vdd _0962_ _0960_ _0947_ _0961_ _0954_ _0955_ vss vdd sky130_fd_sc_hd__a32o_1
XFILLER_24_166 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_62_228 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_47_269 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_46_85 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_46_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_15_100 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_169 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_8 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_7_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_11_361 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2221_ vss vdd d5.fll_core.counter1.count\[9\] _0234_ _0010_ clknet_1_1__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_2
X_2152_ vss vdd d2.t_load\[41\] _0168_ _0402_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_38_225 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1103_ vss vdd _0405_ _0861_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_38_269 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2083_ vss vdd d2.r_reg\[78\] _0099_ _0333_ clknet_4_1_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1034_ vss vdd _0437_ _0824_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1867_ vdd vss _0786_ _0135_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1936_ vdd vss _0792_ _0198_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_21_158 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_21_169 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1798_ vdd vss _0779_ _0073_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_29_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_12_114 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_32_65 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_4_357 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_57_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_35_206 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1721_ vss vdd _0762_ _0013_ _0761_ vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_11_191 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1583_ vss vdd _0662_ d2.r_reg\[23\] _0679_ _0680_ vss vdd sky130_fd_sc_hd__mux2_1
X_1652_ vss vdd _0802_ d2.r_reg\[1\] _0726_ _0727_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_66_342 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2135_ vss vdd d2.t_load\[24\] _0151_ _0385_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2204_ vss vdd d2.t_load\[93\] _0220_ _0454_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2066_ vss vdd d2.r_reg\[61\] _0082_ _0316_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1017_ vss vdd _0814_ d2.r_reg\[84\] net35 _0816_ vss vdd sky130_fd_sc_hd__mux2_1
X_1919_ vdd vss _0791_ _0182_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_1_349 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_1_305 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_57_342 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_27_32 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_17_217 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_40_253 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_40_220 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xclkbuf_4_10_0_clk_in vss vdd clknet_4_10_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
XFILLER_48_342 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_0_382 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1704_ vss vdd _0751_ _0754_ d5.fll_core.counter1.count\[3\] vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_31_264 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1566_ vss vdd _0652_ d2.t_load\[28\] d2.r_reg\[29\] _0668_ vss vdd sky130_fd_sc_hd__mux2_1
X_1497_ vss vdd _0618_ d2.r_reg\[50\] _0620_ _0621_ vss vdd sky130_fd_sc_hd__mux2_1
X_1635_ vss vdd _0262_ _0715_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_54_356 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2049_ vss vdd d2.r_reg\[44\] _0065_ _0299_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2118_ vss vdd d2.t_load\[7\] _0134_ _0368_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_14_209 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_22_253 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_13_89 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_45_301 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_54_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1351_ vss vdd _0520_ _0519_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1420_ vss vdd _0552_ d2.r_reg\[74\] _0567_ _0568_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_63_120 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_304 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1282_ vdd vss _0461_ _0000_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_51_326 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1618_ vss vdd _0684_ d2.r_reg\[12\] _0703_ _0704_ vss vdd sky130_fd_sc_hd__mux2_1
X_0997_ vss vdd _0455_ _0805_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1549_ vss vdd _0289_ _0656_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_39_161 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_10_245 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_10_278 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_65_40 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_46_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1334_ vss vdd _0491_ d5.fll_core.tmp\[4\] _0507_ _0508_ vss vdd sky130_fd_sc_hd__mux2_1
X_1265_ vdd vss d5.fll_core.counter2.count\[1\] _0977_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1403_ vss vdd _0542_ net30 d2.r_reg\[80\] _0556_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_5_293 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_123 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_197 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_120 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xinput3 vss vdd net3 reset vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1196_ vss vdd _0361_ _0910_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_35_76 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_15_326 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_97 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_241 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1050_ vss vdd _0825_ d2.r_reg\[68\] net19 _0833_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_18_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1883_ vdd vss _0787_ _0150_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1952_ vdd vss _0794_ _0212_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1248_ vss vdd d5.fll_core.tmp\[3\] _0961_ d5.fll_core.tmp\[2\] vss vdd sky130_fd_sc_hd__or2_1
X_1317_ vss vdd _0359_ _0494_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XPHY_129 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_118 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_107 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1179_ vss vdd _0369_ _0901_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_24_178 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_24_156 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_270 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XPHY_9 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_62_85 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_62_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_30_159 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_7_69 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2220_ vss vdd d5.fll_core.counter1.count\[8\] _0233_ _0009_ clknet_1_1__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2151_ vss vdd d2.t_load\[40\] _0167_ _0401_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1102_ vss vdd _0859_ d2.r_reg\[44\] d2.t_load\[44\] _0861_ vss vdd sky130_fd_sc_hd__mux2_1
X_2082_ vss vdd d2.r_reg\[77\] _0098_ _0332_ clknet_4_0_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1033_ vss vdd _0814_ d2.r_reg\[76\] net27 _0824_ vss vdd sky130_fd_sc_hd__mux2_1
X_1797_ vdd vss _0779_ _0072_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1866_ vdd vss _0786_ _0134_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1935_ vdd vss _0792_ _0197_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_29_204 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xclkbuf_4_8_0_clk_in vss vdd clknet_4_8_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
XFILLER_4_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1720_ vdd vss d5.fll_core.counter2.count\[0\] d5.fll_core.counter2.count\[2\] _0762_
+ d5.fll_core.counter2.count\[1\] vss vdd sky130_fd_sc_hd__a21oi_1
XFILLER_7_152 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_7_174 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1651_ vss vdd _0519_ d2.t_load\[1\] d2.r_reg\[2\] _0726_ vss vdd sky130_fd_sc_hd__mux2_1
X_1582_ vss vdd _0674_ d2.t_load\[23\] d2.r_reg\[24\] _0679_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_66_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2134_ vss vdd d2.t_load\[23\] _0150_ _0384_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2065_ vss vdd d2.r_reg\[60\] _0081_ _0315_ clknet_4_8_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2203_ vss vdd net43 _0219_ _0453_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1016_ vss vdd _0446_ _0815_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1849_ vdd vss _0784_ _0119_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1918_ vdd vss _0791_ _0181_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_1_317 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_40_210 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_27_44 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_25_273 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_40_232 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_63_324 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_0_361 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_31_221 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_16_240 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_16_295 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1703_ vdd vss _0753_ _0751_ d5.fll_core.counter1.count\[3\] vss vdd sky130_fd_sc_hd__and2_1$1
X_1634_ vss vdd _0706_ d2.r_reg\[7\] _0714_ _0715_ vss vdd sky130_fd_sc_hd__mux2_1
X_1565_ vss vdd _0284_ _0667_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_39_332 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1496_ vss vdd _0608_ d2.t_load\[50\] d2.r_reg\[51\] _0620_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_54_324 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2048_ vss vdd d2.r_reg\[43\] _0064_ _0298_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_39_365 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2117_ vss vdd d2.t_load\[6\] _0133_ _0367_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_13_57 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_49_118 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_1_169 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_54_53 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_54_20 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_45_346 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_225 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1281_ vss vdd _0983_ _0460_ _0461_ _0990_ vss vdd sky130_fd_sc_hd__or3b_1
X_1350_ vss vdd _0519_ net2 vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_0996_ vss vdd _0803_ d2.r_reg\[94\] d2.t_load\[94\] _0805_ vss vdd sky130_fd_sc_hd__mux2_1
X_1617_ vss vdd _0696_ d2.t_load\[12\] d2.r_reg\[13\] _0703_ vss vdd sky130_fd_sc_hd__mux2_1
X_1548_ vss vdd _0640_ d2.r_reg\[34\] _0655_ _0656_ vss vdd sky130_fd_sc_hd__mux2_1
X_1479_ vdd vss _0608_ net2 vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_42_305 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_45_176 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_45_165 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_60_124 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_371 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_5_261 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1402_ vss vdd _0335_ _0555_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1333_ vdd vss _0507_ _0506_ _0502_ vss vdd sky130_fd_sc_hd__and2_1$1
XFILLER_39_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1264_ vdd vss _0976_ _0973_ d2.t_load\[0\] d2.t_load\[5\] _0011_ _0975_ vss vdd
+ sky130_fd_sc_hd__a221o_1
Xinput4 vss vdd net4 s_in vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_51_157 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_51_113 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_24_338 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1195_ vss vdd _0904_ net16 d2.t_load\[0\] _0910_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_35_99 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_35_88 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_27_198 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_33_135 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_21_319 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1882_ vdd vss _0787_ _0149_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1951_ vdd vss _0794_ _0211_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_14_360 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_56_249 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1247_ vss vdd _0959_ _0960_ _0958_ _0956_ vss vdd sky130_fd_sc_hd__o21ai_2
X_1316_ vss vdd _0491_ d5.fll_core.tmp\[8\] _0493_ _0494_ vss vdd sky130_fd_sc_hd__mux2_1
X_1178_ vss vdd _0893_ d2.r_reg\[8\] d2.t_load\[8\] _0901_ vss vdd sky130_fd_sc_hd__mux2_1
XPHY_119 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_108 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_21_57 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_15_113 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_62_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_7_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_7_323 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2150_ vss vdd d2.t_load\[39\] _0166_ _0400_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1101_ vss vdd _0406_ _0860_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1032_ vss vdd _0438_ _0823_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2081_ vss vdd d2.r_reg\[76\] _0097_ _0331_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_61_252 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_61_230 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1934_ vdd vss _0792_ _0196_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_21_105 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1796_ vdd vss _0779_ _0071_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1865_ vdd vss _0786_ _0133_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_16_68 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_8_109 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_20_193 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_35_219 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_43_263 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_28_271 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1581_ vss vdd _0279_ _0678_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_7_186 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1650_ vss vdd _0257_ _0725_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2202_ vss vdd net42 _0218_ _0452_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_21_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_66_377 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2133_ vss vdd d2.t_load\[22\] _0149_ _0383_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2064_ vss vdd d2.r_reg\[59\] _0080_ _0314_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_219 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1015_ vss vdd _0814_ d2.r_reg\[85\] net36 _0815_ vss vdd sky130_fd_sc_hd__mux2_1
X_1917_ vdd vss _0791_ _0772_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1779_ vdd vss _0777_ _0056_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1848_ vdd vss _0784_ _0118_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_1_329 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_48_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_31_277 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1564_ vss vdd _0662_ d2.r_reg\[29\] _0666_ _0667_ vss vdd sky130_fd_sc_hd__mux2_1
X_1702_ vss vdd _0752_ _0003_ _0751_ vss vdd sky130_fd_sc_hd__nor2_1
X_1633_ vss vdd _0696_ d2.t_load\[7\] d2.r_reg\[8\] _0714_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_66_141 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1495_ vss vdd _0306_ _0619_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2047_ vss vdd d2.r_reg\[42\] _0063_ _0297_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2116_ vss vdd d2.t_load\[5\] _0132_ _0366_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_57_196 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_57_141 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_45_369 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_60_317 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_9_237 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_48_152 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1280_ vss vdd _0011_ _0460_ d5.fll_core.counter2.count\[8\] _0991_ d2.t_load\[0\]
+ _0972_ vss vdd sky130_fd_sc_hd__o221a_1
XFILLER_36_358 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_0995_ vss vdd _0456_ _0804_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1547_ vss vdd _0652_ d2.t_load\[34\] d2.r_reg\[35\] _0655_ vss vdd sky130_fd_sc_hd__mux2_1
X_1616_ vss vdd _0268_ _0702_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_5_81 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_39_174 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1478_ vss vdd _0311_ _0607_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_27_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_54_166 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_65_20 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_33_317 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_314 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1401_ vss vdd _0552_ d2.r_reg\[80\] _0554_ _0555_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_5_273 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1332_ vss vdd _0962_ _0506_ _0964_ vss vdd sky130_fd_sc_hd__or2_1
XFILLER_36_133 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1263_ vss vdd d5.fll_core.counter2.count\[3\] _0975_ _0974_ vss vdd sky130_fd_sc_hd__nor2_1
X_1194_ vss vdd _0362_ _0909_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_51_136 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_10_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_269 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_59_225 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_19_79 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_30_309 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_23_383 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1950_ vdd vss _0794_ _0772_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1881_ vdd vss _0787_ _0148_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_51_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1315_ vdd vss _0968_ _0493_ _0950_ vss vdd sky130_fd_sc_hd__xor2_1$1
X_1246_ vdd vss _0943_ _0940_ _0957_ _0959_ vss vdd sky130_fd_sc_hd__a21o_1
X_1177_ vss vdd _0370_ _0900_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_24_103 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XPHY_109 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_20_331 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_250 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_15_169 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_7_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_11_320 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1100_ vss vdd _0859_ d2.r_reg\[45\] d2.t_load\[45\] _0860_ vss vdd sky130_fd_sc_hd__mux2_1
X_1031_ vss vdd _0814_ d2.r_reg\[77\] net28 _0823_ vss vdd sky130_fd_sc_hd__mux2_1
X_2080_ vss vdd d2.r_reg\[75\] _0096_ _0330_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_61_297 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1933_ vdd vss _0792_ _0195_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_21_139 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1795_ vdd vss _0779_ _0773_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1864_ vdd vss _0786_ _0132_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1229_ vss vdd _0926_ _0941_ _0001_ d2.t_load\[20\] _0942_ vss vdd sky130_fd_sc_hd__o211a_1
XFILLER_52_264 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_209 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_12_128 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_20_161 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_4_338 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_11_150 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1580_ vss vdd _0662_ d2.r_reg\[24\] _0677_ _0678_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_7_165 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_7_198 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_66_323 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2132_ vss vdd d2.t_load\[21\] _0148_ _0382_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_14_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2201_ vss vdd net41 _0217_ _0451_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2063_ vss vdd d2.r_reg\[58\] _0079_ _0313_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_34_264 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1014_ vdd vss _0814_ _0802_ vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_19_272 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1847_ vdd vss _0784_ _0117_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1916_ vdd vss _0790_ _0180_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1778_ vdd vss _0777_ _0055_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_57_323 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_27_79 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_25_286 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_63_359 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_48_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_264 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1701_ vdd vss d5.fll_core.counter1.count\[1\] d5.fll_core.counter1.count\[2\] _0752_
+ d5.fll_core.counter1.count\[0\] vss vdd sky130_fd_sc_hd__a21oi_1
X_1563_ vss vdd _0652_ d2.t_load\[29\] d2.r_reg\[30\] _0666_ vss vdd sky130_fd_sc_hd__mux2_1
X_1494_ vss vdd _0618_ d2.r_reg\[51\] _0617_ _0619_ vss vdd sky130_fd_sc_hd__mux2_1
X_1632_ vss vdd _0263_ _0713_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_66_131 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2115_ vss vdd d2.t_load\[4\] _0131_ _0365_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2046_ vss vdd d2.r_reg\[41\] _0062_ _0296_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_22_245 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_49_109 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_57_153 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_38_56 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_205 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_9_249 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_13_267 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_0_193 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_63_134 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_197 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_8_293 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_0994_ vss vdd _0803_ d2.r_reg\[95\] d2.t_load\[95\] _0804_ vss vdd sky130_fd_sc_hd__mux2_1
X_1546_ vss vdd _0290_ _0654_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1615_ vss vdd _0684_ d2.r_reg\[13\] _0701_ _0702_ vss vdd sky130_fd_sc_hd__mux2_1
X_1477_ vss vdd _0596_ d2.r_reg\[56\] _0606_ _0607_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_5_93 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_27_359 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2029_ vss vdd d2.r_reg\[24\] _0045_ _0279_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_65_32 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_45_101 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_65_87 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_26_381 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_60_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1331_ vss vdd _0356_ _0505_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1400_ vss vdd _0542_ net31 d2.r_reg\[81\] _0554_ vss vdd sky130_fd_sc_hd__mux2_1
X_1193_ vss vdd _0904_ d2.r_reg\[1\] d2.t_load\[1\] _0909_ vss vdd sky130_fd_sc_hd__mux2_1
X_1262_ vdd vss d2.t_load\[3\] _0974_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1529_ vss vdd _0640_ d2.r_reg\[40\] _0642_ _0643_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_42_137 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_35_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_23_351 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_65_218 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_18_112 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1880_ vdd vss _0787_ _0147_ vss vdd sky130_fd_sc_hd__inv_2$1
XPHY_90 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_25_90 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_44_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1314_ vss vdd _0360_ _0492_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1245_ vss vdd _0958_ _0940_ _0957_ _0943_ vss vdd sky130_fd_sc_hd__and3_1
XFILLER_49_281 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1176_ vss vdd _0893_ d2.r_reg\[9\] d2.t_load\[9\] _0900_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_20_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_21_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_218 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_30_107 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_23_181 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_7_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xclkbuf_4_13_0_clk_in vss vdd clknet_4_13_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
X_1030_ vss vdd _0439_ _0822_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1932_ vdd vss _0792_ _0194_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1863_ vdd vss _0786_ _0131_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1794_ vdd vss _0778_ _0070_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1228_ vss vdd _0941_ _0917_ _0919_ _0918_ vss vdd sky130_fd_sc_hd__and3_1
XFILLER_29_218 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1159_ vss vdd _0378_ _0890_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_12_107 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_173 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_28_295 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_43_276 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_3_361 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_66_302 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2131_ vss vdd d2.t_load\[20\] _0147_ _0381_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2062_ vss vdd d2.r_reg\[57\] _0078_ _0312_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2200_ vss vdd net40 _0216_ _0450_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_34_221 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1013_ vss vdd _0447_ _0813_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_19_262 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1777_ vdd vss _0777_ _0054_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1915_ vdd vss _0790_ _0179_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1846_ vdd vss _0784_ _0116_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_25_232 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_43_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_4_103 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_48_357 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_16_221 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1700_ vss vdd _0751_ d5.fll_core.counter1.count\[1\] d5.fll_core.counter1.count\[2\]
+ d5.fll_core.counter1.count\[0\] vss vdd sky130_fd_sc_hd__and3_1
X_1631_ vss vdd _0706_ d2.r_reg\[8\] _0712_ _0713_ vss vdd sky130_fd_sc_hd__mux2_1
X_1562_ vss vdd _0285_ _0665_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1493_ vss vdd _0618_ _0892_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_54_349 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2045_ vss vdd d2.r_reg\[40\] _0061_ _0295_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_39_357 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_39_346 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2114_ vss vdd d2.t_load\[3\] _0130_ _0364_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_22_279 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1829_ vdd vss _0783_ _0780_ vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_45_327 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_38_390 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_217 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_21_290 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
Xclkbuf_4_1_0_clk_in vss vdd clknet_4_1_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
XFILLER_63_113 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_0993_ vss vdd _0803_ _0802_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1614_ vss vdd _0696_ d2.t_load\[13\] d2.r_reg\[14\] _0701_ vss vdd sky130_fd_sc_hd__mux2_1
X_1545_ vss vdd _0640_ d2.r_reg\[35\] _0653_ _0654_ vss vdd sky130_fd_sc_hd__mux2_1
X_1476_ vss vdd _0586_ d2.t_load\[56\] d2.r_reg\[57\] _0606_ vss vdd sky130_fd_sc_hd__mux2_1
X_2028_ vss vdd d2.r_reg\[23\] _0044_ _0278_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_39_198 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_35_360 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_24_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_50_341 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_6_209 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_40_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_45_124 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_41_330 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1330_ vss vdd _0491_ d5.fll_core.tmp\[5\] _0504_ _0505_ vss vdd sky130_fd_sc_hd__mux2_1
X_1261_ vdd vss d5.fll_core.counter2.count\[5\] _0973_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1192_ vss vdd _0363_ _0908_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_59_249 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1528_ vss vdd _0630_ d2.t_load\[40\] d2.r_reg\[41\] _0642_ vss vdd sky130_fd_sc_hd__mux2_1
X_1459_ vss vdd _0317_ _0594_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_27_124 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_19_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_42_105 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_35_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_57 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_18_146 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XPHY_91 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_80 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_14_330 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_56_219 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1244_ vdd vss d5.fll_core.tmp\[1\] _0957_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_37_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1313_ vss vdd _0491_ d5.fll_core.tmp\[9\] _0971_ _0492_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_64_296 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1175_ vss vdd _0371_ _0899_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_24_149 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_20_355 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_20_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_21_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_263 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_230 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_296 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_23_193 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_7_337 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1793_ vdd vss _0778_ _0069_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1862_ vdd vss _0786_ _0780_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1931_ vdd vss _0792_ _0193_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1227_ vdd vss d5.fll_core.counter1.count\[0\] _0001_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1158_ vss vdd _0881_ d2.r_reg\[17\] d2.t_load\[17\] _0890_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_37_230 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1089_ vss vdd _0848_ d2.r_reg\[50\] d2.t_load\[50\] _0854_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_32_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_185 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_7_134 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_3_373 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2130_ vss vdd d2.t_load\[19\] _0146_ _0380_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2061_ vss vdd d2.r_reg\[56\] _0077_ _0311_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1012_ vss vdd _0803_ d2.r_reg\[86\] net37 _0813_ vss vdd sky130_fd_sc_hd__mux2_1
X_1914_ vdd vss _0790_ _0178_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_34_277 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_34_244 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1776_ vdd vss _0777_ _0053_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1845_ vdd vss _0784_ _0115_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_25_211 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xclkbuf_1_0__f_vco_in vss vdd clknet_1_0__leaf_vco_in clknet_0_vco_in vss vdd sky130_fd_sc_hd__clkbuf_16
XFILLER_43_69 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_40_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_63_317 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_63_306 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_31_225 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_16_233 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1630_ vss vdd _0696_ d2.t_load\[8\] d2.r_reg\[9\] _0712_ vss vdd sky130_fd_sc_hd__mux2_1
X_1561_ vss vdd _0662_ d2.r_reg\[30\] _0664_ _0665_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_39_303 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1492_ vss vdd _0608_ d2.t_load\[51\] d2.r_reg\[52\] _0617_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_66_177 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_66_155 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2044_ vss vdd d2.r_reg\[39\] _0060_ _0294_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_54_317 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2113_ vss vdd d2.t_load\[2\] _0129_ _0363_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1759_ vdd vss _0775_ _0038_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_1_118 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1828_ vdd vss _0782_ _0100_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_38_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_13_225 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_63_169 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_63_158 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_63_103 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_166 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_0992_ vdd vss _0802_ net1 vss vdd sky130_fd_sc_hd__buf_4$1
X_1544_ vss vdd _0652_ d2.t_load\[35\] d2.r_reg\[36\] _0653_ vss vdd sky130_fd_sc_hd__mux2_1
X_1613_ vss vdd _0269_ _0700_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_5_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1475_ vss vdd _0312_ _0605_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2027_ vss vdd d2.r_reg\[22\] _0043_ _0277_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_54_114 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_49_79 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_45_169 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_60_117 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_386 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_26_372 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_5_221 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1260_ vdd vss d5.fll_core.counter2.count\[0\] _0011_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1191_ vss vdd _0904_ d2.r_reg\[2\] d2.t_load\[2\] _0908_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_36_114 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1527_ vss vdd _0296_ _0641_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_10_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_35_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1458_ vss vdd _0574_ d2.r_reg\[62\] _0593_ _0594_ vss vdd sky130_fd_sc_hd__mux2_1
X_1389_ vss vdd _0339_ _0546_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_19_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_26_191 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_14_320 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_136 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_158 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XPHY_92 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_81 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_70 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_14_353 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1243_ vdd vss d5.fll_core.tmp\[0\] _0956_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1312_ vss vdd _0491_ _0000_ _0483_ _0490_ vss vdd sky130_fd_sc_hd__nand3_4
X_1174_ vss vdd _0893_ d2.r_reg\[10\] d2.t_load\[10\] _0899_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_2_85 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_2_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_64_253 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_32_161 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_21_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_286 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_38_209 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_61_212 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_253 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1930_ vdd vss _0792_ _0192_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1792_ vdd vss _0778_ _0068_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1861_ vdd vss _0785_ _0130_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1226_ vss vdd _0926_ _0939_ _0921_ _0936_ _0940_ vss vdd sky130_fd_sc_hd__a31o_1
X_1157_ vss vdd _0379_ _0889_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_37_275 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_52_278 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_52_245 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1088_ vss vdd _0412_ _0853_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_20_120 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_20_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_57_57 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_7_113 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_3_385 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_34_234 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2060_ vss vdd d2.r_reg\[55\] _0076_ _0310_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1011_ vss vdd _0448_ _0812_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_19_231 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_19_286 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_19_297 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1913_ vdd vss _0790_ _0177_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1775_ vdd vss _0777_ _0052_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1844_ vdd vss _0784_ _0114_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1209_ vss vdd d2.t_load\[29\] d5.fll_core.counter1.count\[9\] _0923_ vss vdd sky130_fd_sc_hd__or2b_1
XFILLER_43_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2189_ vss vdd net29 _0205_ _0439_ clknet_4_1_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_4_116 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_304 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_31_248 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_17_82 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1560_ vss vdd _0652_ d2.t_load\[30\] d2.r_reg\[31\] _0664_ vss vdd sky130_fd_sc_hd__mux2_1
X_1491_ vss vdd _0307_ _0616_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_12_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2112_ vss vdd d2.t_load\[1\] _0128_ _0362_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2043_ vss vdd d2.r_reg\[38\] _0059_ _0293_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1827_ vdd vss _0782_ _0099_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1689_ vss vdd d2.t_load\[44\] d2.t_load\[37\] d2.t_load\[59\] _0746_ vss vdd sky130_fd_sc_hd__mux2_1
X_1758_ vdd vss _0775_ _0037_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_38_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_54_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_13_248 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_21_281 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_0_141 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_0_152 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_351 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_318 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1543_ vss vdd _0652_ net2 vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1612_ vss vdd _0684_ d2.r_reg\[14\] _0699_ _0700_ vss vdd sky130_fd_sc_hd__mux2_1
X_1474_ vss vdd _0596_ d2.r_reg\[57\] _0604_ _0605_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_62_181 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2026_ vss vdd d2.r_reg\[21\] _0042_ _0276_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_50_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_6_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_65_79 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_65_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_65_46 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_26_351 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1190_ vss vdd _0364_ _0907_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_55_90 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_32_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_32_332 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1526_ vss vdd _0640_ d2.r_reg\[41\] _0639_ _0641_ vss vdd sky130_fd_sc_hd__mux2_1
X_1457_ vss vdd _0586_ d2.t_load\[62\] d2.r_reg\[63\] _0593_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_35_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_27_137 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1388_ vss vdd _0530_ d2.r_reg\[84\] _0545_ _0546_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_19_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_51_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_42_129 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_23_376 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2009_ vss vdd d2.r_reg\[4\] _0025_ _0259_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_2_258 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XPHY_82 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_71 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_60 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_14_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XPHY_93 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_184 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_41_151 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1311_ vss vdd _0490_ _0482_ _0489_ _0946_ _0485_ vss vdd sky130_fd_sc_hd__o31a_1
XFILLER_49_240 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1242_ vss vdd _0945_ _0955_ d5.fll_core.tmp\[2\] vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1173_ vss vdd _0372_ _0898_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_2_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_17_181 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_302 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1509_ vss vdd _0618_ d2.r_reg\[46\] _0628_ _0629_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_46_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_15_107 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_62_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_11_368 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_36_92 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_70 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1860_ vdd vss _0785_ _0129_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_52_91 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1791_ vdd vss _0778_ _0067_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_42_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1225_ vss vdd _0934_ _0937_ _0931_ _0939_ _0938_ _0926_ vss vdd sky130_fd_sc_hd__a41o_1
X_1156_ vss vdd _0881_ d2.r_reg\[18\] d2.t_load\[18\] _0889_ vss vdd sky130_fd_sc_hd__mux2_1
X_1087_ vss vdd _0848_ d2.r_reg\[51\] d2.t_load\[51\] _0853_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_16_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1989_ vdd vss _0801_ _0239_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_57_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_28_221 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_11_121 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_11_165 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_22_50 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_66_316 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_66_349 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1010_ vss vdd _0803_ d2.r_reg\[87\] net38 _0812_ vss vdd sky130_fd_sc_hd__mux2_1
X_1912_ vdd vss _0790_ _0176_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_8_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_8_85 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1843_ vdd vss _0784_ _0113_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1774_ vdd vss _0777_ _0051_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_6_180 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1208_ vss vdd d2.t_load\[28\] d5.fll_core.counter1.count\[8\] _0922_ vss vdd sky130_fd_sc_hd__or2b_1
XFILLER_57_349 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1139_ vss vdd _0870_ d2.r_reg\[26\] d2.t_load\[26\] _0880_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_43_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2188_ vss vdd net28 _0204_ _0438_ clknet_4_1_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_33_71 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_31_205 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1490_ vss vdd _0596_ d2.r_reg\[52\] _0615_ _0616_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_66_124 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_66_113 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2042_ vss vdd d2.r_reg\[37\] _0058_ _0292_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_3_194 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2111_ vss vdd d2.t_load\[0\] _0127_ _0361_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_47_360 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_22_238 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_282 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1826_ vdd vss _0782_ _0098_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1688_ vss vdd net10 _0745_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1757_ vdd vss _0775_ _0036_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_57_113 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_45_308 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_13_205 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_0_186 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_60_80 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1611_ vss vdd _0696_ d2.t_load\[14\] d2.r_reg\[15\] _0699_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_8_253 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1542_ vss vdd _0291_ _0651_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1473_ vss vdd _0586_ d2.t_load\[57\] d2.r_reg\[58\] _0604_ vss vdd sky130_fd_sc_hd__mux2_1
X_2025_ vss vdd d2.r_reg\[20\] _0041_ _0275_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_39_113 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_50_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_24_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1809_ vdd vss _0781_ _0082_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_49_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_65_69 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_53_160 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_5_201 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_32_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_219 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1525_ vss vdd _0640_ _0892_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1456_ vss vdd _0318_ _0592_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1387_ vss vdd _0542_ net35 d2.r_reg\[85\] _0545_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_35_182 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_35_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_27_105 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2008_ vss vdd d2.r_reg\[3\] _0024_ _0258_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_51_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_23_344 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_248 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_105 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_94 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_83 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_72 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_61 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_50 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_14_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1241_ vss vdd _0945_ _0954_ d5.fll_core.tmp\[3\] vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1310_ vss vdd _0489_ d5.fll_core.tmp\[3\] _0488_ _0946_ vss vdd sky130_fd_sc_hd__nand3_1
XFILLER_1_281 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1172_ vss vdd _0893_ d2.r_reg\[11\] d2.t_load\[11\] _0898_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_2_98 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_65 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_32_185 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_32_152 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_17_193 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1508_ vss vdd _0608_ d2.t_load\[46\] d2.r_reg\[47\] _0628_ vss vdd sky130_fd_sc_hd__mux2_1
X_1439_ vss vdd _0574_ d2.r_reg\[68\] _0580_ _0581_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_62_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_277 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_2_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_46_222 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1790_ vdd vss _0778_ _0066_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_14_141 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_14_130 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1224_ vdd vss _0938_ _0922_ _0924_ _0923_ vss vdd sky130_fd_sc_hd__a21boi_1
XFILLER_35_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1155_ vss vdd _0380_ _0888_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_37_255 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1086_ vss vdd _0413_ _0852_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_32_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1988_ vdd vss _0801_ _0238_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_57_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_43_225 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
Xclkbuf_4_4_0_clk_in vss vdd clknet_4_4_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
X_1773_ vdd vss _0777_ _0773_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1911_ vdd vss _0790_ _0175_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_8_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_8_97 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1842_ vdd vss _0784_ _0112_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_6_192 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1207_ vss vdd _0914_ _0916_ _0921_ _0913_ _0920_ vss vdd sky130_fd_sc_hd__o22ai_1
X_2187_ vss vdd net27 _0203_ _0437_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_2
X_1138_ vss vdd _0388_ _0879_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_43_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1069_ vss vdd _0836_ d2.r_reg\[59\] d2.t_load\[59\] _0843_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_25_247 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_25_225 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_129 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_17_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_17_95 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_66_169 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_66_103 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2041_ vss vdd d2.r_reg\[36\] _0057_ _0291_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2110_ vss vdd d5.fll_core.tmp\[9\] _0126_ _0360_ clknet_1_0__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfrtp_2
X_1756_ vdd vss _0775_ _0035_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1825_ vdd vss _0782_ _0097_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1687_ vss vdd d2.t_load\[44\] d2.t_load\[36\] d2.t_load\[58\] _0745_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_65_191 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_57_169 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2239_ vss vdd d2.t_load\[63\] _0252_ d5.mux01.out\[7\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
XFILLER_13_217 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_21_250 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_48_103 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_29_350 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_28_94 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1610_ vss vdd _0270_ _0698_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_8_221 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_8_265 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1541_ vss vdd _0640_ d2.r_reg\[36\] _0650_ _0651_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_39_125 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1472_ vss vdd _0313_ _0603_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2024_ vss vdd d2.r_reg\[19\] _0040_ _0274_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_47_180 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_50_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_50_334 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_10_209 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_49_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_40_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1808_ vdd vss _0781_ _0081_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1739_ vss vdd _0773_ _0772_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_60_109 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_323 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_213 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_14_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_14_74 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_106 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_29_191 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_17_320 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_17_342 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_32_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1524_ vss vdd _0630_ d2.t_load\[41\] d2.r_reg\[42\] _0639_ vss vdd sky130_fd_sc_hd__mux2_1
X_1455_ vss vdd _0574_ d2.r_reg\[63\] _0591_ _0592_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_4_290 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1386_ vss vdd _0340_ _0544_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_35_150 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2007_ vss vdd d2.r_reg\[2\] _0023_ _0257_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_51_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_2_205 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_58_297 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_58_253 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XPHY_95 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_84 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_73 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_62 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_51 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_25_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_14_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_40 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_49_253 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1171_ vss vdd _0373_ _0897_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1240_ vdd vss _0953_ _0952_ _0951_ vss vdd sky130_fd_sc_hd__and2_1$1
XFILLER_2_77 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_1_293 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1507_ vss vdd _0302_ _0627_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_55_212 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1369_ vss vdd _0530_ d2.r_reg\[90\] _0532_ _0533_ vss vdd sky130_fd_sc_hd__mux2_1
X_1438_ vss vdd _0564_ net19 d2.r_reg\[69\] _0580_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_11_348 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_245 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_10_370 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_14_153 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_14_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1223_ vss vdd _0937_ _0933_ _0928_ _0932_ _0929_ vss vdd sky130_fd_sc_hd__a211o_1
X_1154_ vss vdd _0881_ d2.r_reg\[19\] d2.t_load\[19\] _0888_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_28_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1085_ vss vdd _0848_ d2.r_reg\[52\] d2.t_load\[52\] _0852_ vss vdd sky130_fd_sc_hd__mux2_1
X_1987_ vdd vss _0801_ _0237_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_57_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_43_248 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_51_292 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_51_281 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_7_105 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_22_41 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_22_74 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_22_85 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_63_81 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1910_ vdd vss _0790_ _0174_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1772_ vdd vss _0776_ _0050_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_8_65 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1841_ vdd vss _0784_ _0111_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1137_ vss vdd _0870_ d2.r_reg\[27\] d2.t_load\[27\] _0879_ vss vdd sky130_fd_sc_hd__mux2_1
X_1206_ vdd vss _0920_ _0917_ _0919_ _0918_ vss vdd sky130_fd_sc_hd__a21boi_1
XFILLER_25_204 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2186_ vss vdd net26 _0202_ _0436_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1068_ vss vdd _0421_ _0842_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_33_292 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_318 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_33_84 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_66_148 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2040_ vss vdd d2.r_reg\[35\] _0056_ _0290_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_62_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1686_ vss vdd net9 _0744_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1755_ vdd vss _0775_ _0034_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1824_ vdd vss _0782_ _0096_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_38_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2238_ vss vdd d2.t_load\[62\] _0251_ d5.mux01.out\[6\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
XFILLER_53_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2169_ vss vdd d2.t_load\[58\] _0185_ _0419_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_56_181 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_159 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_365 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1540_ vss vdd _0630_ d2.t_load\[36\] d2.r_reg\[37\] _0650_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_8_233 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1471_ vss vdd _0596_ d2.r_reg\[58\] _0602_ _0603_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_10_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2023_ vss vdd d2.r_reg\[18\] _0039_ _0273_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_50_357 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1807_ vdd vss _0781_ _0780_ vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_49_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1669_ vss vdd _0847_ d2.t_load\[48\] d5.fll_core.tmp\[3\] _0736_ vss vdd sky130_fd_sc_hd__mux2_1
X_1738_ vdd vss _0772_ net3 vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_38_192 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_74 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_30_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_5_225 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_58_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1523_ vss vdd _0297_ _0638_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1454_ vss vdd _0586_ d2.t_load\[63\] d2.r_reg\[64\] _0591_ vss vdd sky130_fd_sc_hd__mux2_1
X_1385_ vss vdd _0530_ d2.r_reg\[85\] _0543_ _0544_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_35_140 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_23_313 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2006_ vss vdd d2.r_reg\[1\] _0022_ _0256_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_58_232 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_228 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_58_287 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_30 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_96 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_85 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_74 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_63 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_52 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_14_346 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_41 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1170_ vss vdd _0893_ d2.r_reg\[12\] d2.t_load\[12\] _0897_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_1_261 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_64_279 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_17_140 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1506_ vss vdd _0618_ d2.r_reg\[47\] _0626_ _0627_ vss vdd sky130_fd_sc_hd__mux2_1
X_1437_ vss vdd _0324_ _0579_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1299_ vss vdd d2.t_load\[16\] d5.fll_core.counter1.count\[6\] _0478_ _0474_ vss
+ vdd sky130_fd_sc_hd__or3b_1
XFILLER_46_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1368_ vss vdd _0520_ net41 d2.r_reg\[91\] _0532_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_11_327 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_11_87 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_61_238 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_279 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_10_382 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_14_165 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1222_ vss vdd _0936_ _0931_ _0935_ vss vdd sky130_fd_sc_hd__and2b_1
X_1153_ vss vdd _0381_ _0887_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_37_268 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1084_ vss vdd _0414_ _0851_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_52_238 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1986_ vdd vss _0801_ _0236_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_57_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_36_290 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_11_113 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_59_371 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_42_271 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1840_ vss vdd _0784_ _0780_ vss vdd sky130_fd_sc_hd__clkbuf_8
X_1771_ vdd vss _0776_ _0049_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_8_77 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_10_190 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_57_308 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1136_ vss vdd _0389_ _0878_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1205_ vss vdd d2.t_load\[21\] d5.fll_core.counter1.count\[1\] _0919_ vss vdd sky130_fd_sc_hd__or2b_1
X_1067_ vss vdd _0836_ d2.r_reg\[60\] d2.t_load\[60\] _0842_ vss vdd sky130_fd_sc_hd__mux2_1
X_2185_ vss vdd net25 _0201_ _0435_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1969_ vdd vss _0798_ _0796_ d5.fll_core.corner_tmp\[1\] vss vdd sky130_fd_sc_hd__and2_1$1
XFILLER_33_271 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_24_293 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_17_75 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_3_142 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_62_355 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_62_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1823_ vdd vss _0782_ _0095_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1685_ vss vdd d2.t_load\[44\] d2.t_load\[35\] d2.t_load\[57\] _0744_ vss vdd sky130_fd_sc_hd__mux2_1
X_1754_ vdd vss _0775_ _0033_ vss vdd sky130_fd_sc_hd__inv_2$1
X_2237_ vss vdd d2.t_load\[61\] _0250_ d5.mux01.out\[5\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
XFILLER_65_160 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1119_ vss vdd _0397_ _0869_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_54_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_53_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2168_ vss vdd d2.t_load\[57\] _0184_ _0418_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2099_ vss vdd d2.r_reg\[94\] _0115_ _0349_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_48_116 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_28_85 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_28_41 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_8_245 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1470_ vss vdd _0586_ d2.t_load\[58\] d2.r_reg\[59\] _0602_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_39_149 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_62_174 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_62_141 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2022_ vss vdd d2.r_reg\[17\] _0038_ _0272_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_35_311 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1806_ vdd vss _0780_ _0772_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1599_ vss vdd _0684_ d2.r_reg\[18\] _0690_ _0691_ vss vdd sky130_fd_sc_hd__mux2_1
X_1668_ vss vdd d5.mux01.out\[2\] _0735_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1737_ vdd vss _0770_ _0020_ d5.fll_core.counter2.count\[9\] vss vdd sky130_fd_sc_hd__xor2_1$1
XFILLER_38_171 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_26_344 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_26_300 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_53_174 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_358 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_237 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_39_84 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_39_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_83 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_141 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1522_ vss vdd _0618_ d2.r_reg\[42\] _0637_ _0638_ vss vdd sky130_fd_sc_hd__mux2_1
X_1453_ vss vdd _0319_ _0590_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1384_ vss vdd _0542_ net36 d2.r_reg\[86\] _0543_ vss vdd sky130_fd_sc_hd__mux2_1
X_2005_ vss vdd net16 _0021_ _0255_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XPHY_64 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_53 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_26_130 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_20 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_31 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_42 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_97 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_86 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_177 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_75 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_64_236 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_1_273 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_17_152 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1505_ vss vdd _0608_ d2.t_load\[47\] d2.r_reg\[48\] _0626_ vss vdd sky130_fd_sc_hd__mux2_1
X_1436_ vss vdd _0574_ d2.r_reg\[69\] _0578_ _0579_ vss vdd sky130_fd_sc_hd__mux2_1
X_1367_ vss vdd _0346_ _0531_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1298_ vdd vss d5.fll_core.counter1.count\[8\] _0477_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_62_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_36_85 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_14_177 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_6_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1221_ vdd vss _0935_ _0934_ _0933_ _0932_ d5.fll_core.counter1.count\[4\] _0927_
+ vss vdd sky130_fd_sc_hd__o2111a_1
X_1152_ vss vdd _0881_ d2.r_reg\[20\] d2.t_load\[20\] _0887_ vss vdd sky130_fd_sc_hd__mux2_1
X_1083_ vss vdd _0848_ d2.r_reg\[53\] d2.t_load\[53\] _0851_ vss vdd sky130_fd_sc_hd__mux2_1
X_1985_ vdd vss _0801_ _0235_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_9_181 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_28_236 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_28_214 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1419_ vss vdd _0564_ net25 d2.r_reg\[75\] _0567_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_28_258 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_22_98 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_3_324 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_383 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_19_225 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1770_ vdd vss _0776_ _0048_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1204_ vss vdd d5.fll_core.counter1.count\[1\] d2.t_load\[21\] _0918_ vss vdd sky130_fd_sc_hd__or2b_1
X_2184_ vss vdd net24 _0200_ _0434_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1135_ vss vdd _0870_ d2.r_reg\[28\] d2.t_load\[28\] _0878_ vss vdd sky130_fd_sc_hd__mux2_1
X_1066_ vss vdd _0422_ _0841_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1899_ vdd vss _0789_ _0164_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1968_ vss vdd _0457_ _0797_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_0_349 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_0_305 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_56_320 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_33_20 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_180 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_62_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_47_353 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_15_261 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_22_209 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1753_ vdd vss _0775_ _0032_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_30_275 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1822_ vdd vss _0782_ _0094_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1684_ vss vdd net8 _0743_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_57_106 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2236_ vss vdd d2.t_load\[60\] _0249_ d5.mux01.out\[4\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
X_2167_ vss vdd d2.t_load\[56\] _0183_ _0417_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1118_ vss vdd _0859_ d2.r_reg\[36\] d2.t_load\[36\] _0869_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_53_389 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_53_356 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2098_ vss vdd d2.r_reg\[93\] _0114_ _0348_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1049_ vss vdd _0430_ _0832_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_0_135 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_29_375 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_44_85 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_12_253 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_5_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2021_ vss vdd d2.r_reg\[16\] _0037_ _0271_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_62_197 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_50_348 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_35_389 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1805_ vdd vss _0779_ _0080_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1736_ vss vdd _0771_ _0019_ _0770_ vss vdd sky130_fd_sc_hd__nor2_1
X_1598_ vss vdd _0674_ d2.t_load\[18\] d2.r_reg\[19\] _0690_ vss vdd sky130_fd_sc_hd__mux2_1
X_1667_ vss vdd _0847_ d2.t_load\[47\] d5.fll_core.tmp\[2\] _0735_ vss vdd sky130_fd_sc_hd__mux2_1
X_2219_ vss vdd d5.fll_core.counter1.count\[7\] _0232_ _0008_ clknet_1_1__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_334 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_41_337 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_5_249 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_62 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_197 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_17_367 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1521_ vss vdd _0630_ d2.t_load\[42\] d2.r_reg\[43\] _0637_ vss vdd sky130_fd_sc_hd__mux2_1
X_1452_ vss vdd _0574_ d2.r_reg\[64\] _0589_ _0590_ vss vdd sky130_fd_sc_hd__mux2_1
X_1383_ vss vdd _0542_ _0519_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_2004_ vdd vss _0773_ _0254_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1719_ vss vdd _0761_ d5.fll_core.counter2.count\[1\] d5.fll_core.counter2.count\[0\]
+ d5.fll_core.counter2.count\[2\] vss vdd sky130_fd_sc_hd__and3_1
XFILLER_58_245 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XPHY_98 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_87 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_145 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_76 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_65 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_54 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_10 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_21 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_32 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_43 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_97 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xclkbuf_4_7_0_clk_in vss vdd clknet_4_7_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
XFILLER_64_204 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_49_289 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_17_164 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_330 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_63_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1504_ vss vdd _0303_ _0625_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1435_ vss vdd _0564_ net20 d2.r_reg\[70\] _0578_ vss vdd sky130_fd_sc_hd__mux2_1
X_1366_ vss vdd _0530_ d2.r_reg\[91\] _0529_ _0531_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_55_237 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1297_ vss vdd _0476_ _0463_ _0474_ d2.t_load\[15\] _0475_ vss vdd sky130_fd_sc_hd__a211o_1
XFILLER_23_156 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_46_215 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_52_85 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_52_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_14_189 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_6_344 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_6_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1220_ vss vdd d5.fll_core.counter1.count\[7\] d2.t_load\[27\] _0934_ vss vdd sky130_fd_sc_hd__or2b_1
X_1151_ vss vdd _0382_ _0886_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1082_ vss vdd _0415_ _0850_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1984_ vdd vss _0801_ d5.fll_core.counter_reset vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_9_193 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_137 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1349_ vss vdd _0491_ _0351_ d5.fll_core.tmp\[0\] vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1418_ vss vdd _0330_ _0566_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_11_137 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_7_119 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_63_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_6_152 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_65_310 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1134_ vss vdd _0390_ _0877_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1203_ vss vdd d5.fll_core.counter1.count\[0\] d2.t_load\[20\] _0917_ vss vdd sky130_fd_sc_hd__or2b_1
XFILLER_26_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2183_ vss vdd net23 _0199_ _0433_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1065_ vss vdd _0836_ d2.r_reg\[61\] d2.t_load\[61\] _0841_ vss vdd sky130_fd_sc_hd__mux2_1
X_1898_ vdd vss _0789_ _0163_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1967_ vss vdd _0796_ d5.fll_core.corner_tmp\[0\] _0947_ _0797_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_0_317 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_56_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_33_65 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_33_32 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_24_262 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_62_324 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1683_ vss vdd d2.t_load\[44\] d2.t_load\[34\] d2.t_load\[56\] _0743_ vss vdd sky130_fd_sc_hd__mux2_1
X_1752_ vdd vss _0775_ _0031_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1821_ vdd vss _0782_ _0093_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1117_ vss vdd _0398_ _0868_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2235_ vss vdd d2.t_load\[59\] _0248_ d5.mux01.out\[3\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
XFILLER_38_365 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_38_321 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2166_ vss vdd d2.t_load\[55\] _0182_ _0416_ clknet_4_9_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2097_ vss vdd d2.r_reg\[92\] _0113_ _0347_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1048_ vss vdd _0825_ d2.r_reg\[69\] net20 _0832_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_0_103 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_48_129 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_29_343 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_28_54 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_0_169 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_44_75 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_29_387 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_12_221 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_60_96 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_60_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_12_276 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_69 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_151 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2020_ vss vdd d2.r_reg\[15\] _0036_ _0270_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_35_346 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_35_324 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_50_327 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1666_ vss vdd d5.mux01.out\[1\] _0734_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1804_ vdd vss _0779_ _0079_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1735_ vdd vss d5.fll_core.counter2.count\[7\] d5.fll_core.counter2.count\[8\] _0771_
+ _0768_ vss vdd sky130_fd_sc_hd__a21oi_1
X_1597_ vss vdd _0274_ _0689_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2218_ vss vdd d5.fll_core.counter1.count\[6\] _0231_ _0007_ clknet_1_1__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_2
X_2149_ vss vdd d2.t_load\[38\] _0165_ _0399_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_53_187 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_349 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_316 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_39_97 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_154 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_40_360 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_17_379 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1520_ vss vdd _0298_ _0636_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1451_ vss vdd _0586_ d2.t_load\[64\] d2.r_reg\[65\] _0589_ vss vdd sky130_fd_sc_hd__mux2_1
X_1382_ vss vdd _0341_ _0541_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_35_121 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2003_ vdd vss _0773_ _0253_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_23_327 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_50_179 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_50_168 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_31_371 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1718_ vdd vss d5.fll_core.counter2.count\[1\] _0012_ d5.fll_core.counter2.count\[0\]
+ vss vdd sky130_fd_sc_hd__xor2_1$1
X_1649_ vss vdd _0706_ d2.r_reg\[2\] _0724_ _0725_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_58_279 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XPHY_99 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_88 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_124 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_77 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_66 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_55 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_25_77 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_11 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_22 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_14_305 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_33 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_44 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_49_202 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_9_364 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_56_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1503_ vss vdd _0618_ d2.r_reg\[48\] _0624_ _0625_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_55_205 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1296_ vdd vss d5.fll_core.counter1.count\[6\] _0475_ d2.t_load\[16\] vss vdd sky130_fd_sc_hd__xor2_1$1
X_1434_ vss vdd _0325_ _0577_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1365_ vdd vss _0530_ _0892_ vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_48_290 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_11_79 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_61_219 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_46_238 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_52_53 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1150_ vss vdd _0881_ d2.r_reg\[21\] d2.t_load\[21\] _0886_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_37_216 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_52_208 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1081_ vss vdd _0848_ d2.r_reg\[54\] d2.t_load\[54\] _0850_ vss vdd sky130_fd_sc_hd__mux2_1
X_1983_ vdd vss _0800_ _0234_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_20_149 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1417_ vss vdd _0552_ d2.r_reg\[75\] _0565_ _0566_ vss vdd sky130_fd_sc_hd__mux2_1
X_1348_ vss vdd _0352_ _0518_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_28_249 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1279_ vss vdd _0985_ _0991_ d5.fll_core.counter2.count\[4\] d2.t_load\[2\] _0984_
+ vss vdd sky130_fd_sc_hd__o22a_1
XFILLER_51_252 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_3_337 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_3_304 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_47_20 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_86 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_27_260 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_19_249 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_6_131 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_6_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_65_366 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_65_300 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1133_ vss vdd _0870_ d2.r_reg\[29\] d2.t_load\[29\] _0877_ vss vdd sky130_fd_sc_hd__mux2_1
X_1202_ vdd vss _0915_ _0911_ _0916_ _0912_ _0914_ vss vdd sky130_fd_sc_hd__or4_1
X_1064_ vss vdd _0423_ _0840_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2182_ vss vdd net22 _0198_ _0432_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_19_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1966_ vdd vss _0772_ _0796_ _0461_ _0490_ vss vdd sky130_fd_sc_hd__or3_1
X_1897_ vdd vss _0789_ _0162_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_0_329 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_56_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_33_44 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_193 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_58_96 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_58_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_388 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1820_ vdd vss _0782_ _0092_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_15_274 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1751_ vdd vss _0775_ _0773_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1682_ vss vdd d5.mux01.out\[9\] _0742_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_30_299 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2234_ vss vdd d2.t_load\[58\] _0247_ d5.mux01.out\[2\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
X_1116_ vss vdd _0859_ d2.r_reg\[37\] d2.t_load\[37\] _0868_ vss vdd sky130_fd_sc_hd__mux2_1
X_2165_ vss vdd d2.t_load\[54\] _0181_ _0415_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1047_ vss vdd _0431_ _0831_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2096_ vss vdd d2.r_reg\[91\] _0112_ _0346_ clknet_4_7_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1949_ vdd vss _0793_ _0210_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_56_141 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_44_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_0_159 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_336 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_44_65 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_12_233 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_60_53 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_60_20 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_5_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_35_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1803_ vdd vss _0779_ _0078_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1596_ vss vdd _0684_ d2.r_reg\[19\] _0688_ _0689_ vss vdd sky130_fd_sc_hd__mux2_1
X_1665_ vss vdd _0847_ d2.t_load\[46\] d5.fll_core.tmp\[1\] _0734_ vss vdd sky130_fd_sc_hd__mux2_1
X_1734_ vss vdd _0770_ d5.fll_core.counter2.count\[8\] d5.fll_core.counter2.count\[7\]
+ _0768_ vss vdd sky130_fd_sc_hd__and3_1
XFILLER_7_292 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2217_ vss vdd d5.fll_core.counter1.count\[5\] _0230_ _0006_ clknet_1_1__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_38_141 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_2148_ vss vdd d2.t_load\[37\] _0164_ _0398_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_53_133 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_26_358 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2079_ vss vdd d2.r_reg\[74\] _0095_ _0329_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_44_166 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_65_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1450_ vss vdd _0320_ _0588_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1381_ vss vdd _0530_ d2.r_reg\[86\] _0540_ _0541_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_50_103 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2002_ vdd vss _0773_ _0252_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_31_383 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1717_ vdd vss _0759_ _0010_ d5.fll_core.counter1.count\[9\] vss vdd sky130_fd_sc_hd__xor2_1$1
X_1579_ vss vdd _0674_ d2.t_load\[24\] d2.r_reg\[25\] _0677_ vss vdd sky130_fd_sc_hd__mux2_1
X_1648_ vss vdd _0519_ d2.t_load\[2\] d2.r_reg\[3\] _0724_ vss vdd sky130_fd_sc_hd__mux2_1
XPHY_12 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_89 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_158 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_78 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_67 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_56 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_26_166 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_23 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_34 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_22_361 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_45 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_49_225 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_66_96 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_66_85 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_66_74 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_64_228 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_32_125 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_376 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_49_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1502_ vss vdd _0608_ d2.t_load\[48\] d2.r_reg\[49\] _0624_ vss vdd sky130_fd_sc_hd__mux2_1
X_1433_ vss vdd _0574_ d2.r_reg\[70\] _0576_ _0577_ vss vdd sky130_fd_sc_hd__mux2_1
X_1295_ vdd vss _0474_ _0473_ d2.t_load\[17\] vss vdd sky130_fd_sc_hd__and2_1$1
X_1364_ vss vdd _0520_ net42 d2.r_reg\[92\] _0529_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_63_261 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_23_169 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_31_180 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_54_294 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_54_283 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_99 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_77 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_10_320 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_6_357 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1080_ vss vdd _0416_ _0849_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1982_ vdd vss _0800_ _0233_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_60_264 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_162 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1347_ vss vdd _0491_ d5.fll_core.tmp\[1\] _0517_ _0518_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_3_81 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1416_ vss vdd _0564_ net26 d2.r_reg\[76\] _0565_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_36_283 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1278_ vss vdd _0990_ d5.fll_core.counter2.count\[4\] _0988_ _0984_ _0989_ vss vdd
+ sky130_fd_sc_hd__a211o_1
XFILLER_51_275 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_3_349 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_32 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_19_206 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_42_297 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_42_264 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_8_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_10_161 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1201_ vss vdd _0915_ d5.fll_core.counter1.count\[2\] d2.t_load\[22\] vss vdd sky130_fd_sc_hd__and2b_1
XFILLER_65_378 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1132_ vss vdd _0391_ _0876_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1063_ vss vdd _0836_ d2.r_reg\[62\] d2.t_load\[62\] _0840_ vss vdd sky130_fd_sc_hd__mux2_1
X_2181_ vss vdd net21 _0197_ _0431_ clknet_4_0_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1965_ vdd vss _0795_ _0224_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1896_ vdd vss _0789_ _0161_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_56_345 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_56_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_24_286 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_24_253 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_16_209 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_17_68 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_58_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_3_113 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_62_348 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_62_304 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_47_345 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1750_ vdd vss _0774_ _0030_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1681_ vss vdd d2.t_load\[55\] d2.t_load\[54\] d5.fll_core.tmp\[9\] _0742_ vss vdd
+ sky130_fd_sc_hd__mux2_1
X_2233_ vss vdd d2.t_load\[57\] _0246_ d5.mux01.out\[1\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
XFILLER_31_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2164_ vss vdd d2.t_load\[53\] _0180_ _0414_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1115_ vss vdd _0399_ _0867_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_53_348 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_38_356 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1046_ vss vdd _0825_ d2.r_reg\[70\] net21 _0831_ vss vdd sky130_fd_sc_hd__mux2_1
X_2095_ vss vdd d2.r_reg\[90\] _0111_ _0345_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1879_ vdd vss _0787_ _0146_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1948_ vdd vss _0793_ _0209_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_28_78 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_28_67 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_12_245 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_5_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_131 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_62_101 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_50_318 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_47_164 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1802_ vdd vss _0779_ _0077_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1733_ vss vdd _0768_ _0018_ _0980_ vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1595_ vss vdd _0674_ d2.t_load\[19\] d2.r_reg\[20\] _0688_ vss vdd sky130_fd_sc_hd__mux2_1
X_1664_ vss vdd d5.mux01.out\[0\] _0733_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2147_ vss vdd d2.t_load\[36\] _0163_ _0397_ clknet_4_10_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2216_ vss vdd d5.fll_core.counter1.count\[4\] _0229_ _0005_ clknet_1_1__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_38_197 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_38_186 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_38_164 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_307 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1029_ vss vdd _0814_ d2.r_reg\[78\] net29 _0822_ vss vdd sky130_fd_sc_hd__mux2_1
X_2078_ vss vdd d2.r_reg\[73\] _0094_ _0328_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_55_76 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_112 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_241 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1380_ vss vdd _0520_ net37 d2.r_reg\[87\] _0540_ vss vdd sky130_fd_sc_hd__mux2_1
X_2001_ vdd vss _0773_ _0251_ vss vdd sky130_fd_sc_hd__inv_2$1
Xclkbuf_4_12_0_clk_in vss vdd clknet_4_12_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
XFILLER_16_370 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1716_ vss vdd _0760_ _0009_ _0759_ vss vdd sky130_fd_sc_hd__nor2_1
X_1578_ vss vdd _0280_ _0676_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1647_ vss vdd _0258_ _0723_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_66_281 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XPHY_13 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_24 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_35 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_46 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_137 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XPHY_79 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_68 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_57 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_25_68 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_41_89 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_66_42 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_57_281 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_32_104 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_388 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1501_ vss vdd _0304_ _0623_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1432_ vss vdd _0564_ net21 d2.r_reg\[71\] _0576_ vss vdd sky130_fd_sc_hd__mux2_1
X_1363_ vss vdd _0347_ _0528_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1294_ vdd vss d5.fll_core.counter1.count\[7\] _0473_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_11_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_45_262 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1981_ vdd vss _0800_ _0232_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_60_287 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_60_232 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_9_130 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_13_181 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_61_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1346_ vss vdd _0516_ _0517_ _0956_ vss vdd sky130_fd_sc_hd__xnor2_1$1
XFILLER_28_229 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_3_93 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1415_ vss vdd _0564_ _0519_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1277_ vss vdd _0974_ d2.t_load\[5\] _0973_ _0989_ d5.fll_core.counter2.count\[3\]
+ vss vdd sky130_fd_sc_hd__a2bb2o_1
XFILLER_51_265 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_3_317 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_47_44 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_19_218 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_27_273 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1200_ vss vdd _0914_ d5.fll_core.counter1.count\[3\] d2.t_load\[23\] vss vdd sky130_fd_sc_hd__and2b_1
XFILLER_40_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2180_ vss vdd net20 _0196_ _0430_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1131_ vss vdd _0870_ d2.r_reg\[30\] d2.t_load\[30\] _0876_ vss vdd sky130_fd_sc_hd__mux2_1
X_1062_ vss vdd _0424_ _0839_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1895_ vdd vss _0789_ _0780_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1964_ vdd vss _0795_ _0223_ vss vdd sky130_fd_sc_hd__inv_2$1
Xclkbuf_4_0_0_clk_in vss vdd clknet_4_0_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
X_1329_ vdd vss _0503_ _0504_ _0963_ vss vdd sky130_fd_sc_hd__xor2_1$1
XFILLER_33_57 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_24_243 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_58_65 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_3_169 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1680_ vss vdd d5.mux01.out\[8\] _0741_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_65_132 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1114_ vss vdd _0859_ d2.r_reg\[38\] d2.t_load\[38\] _0867_ vss vdd sky130_fd_sc_hd__mux2_1
X_2232_ vss vdd d2.t_load\[56\] _0245_ d5.mux01.out\[0\] d5.fll_core.strobe vss vdd
+ sky130_fd_sc_hd__dfrtp_1$1
X_2163_ vss vdd d2.t_load\[52\] _0179_ _0413_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_24_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_65_198 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_61_371 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1045_ vss vdd _0432_ _0830_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2094_ vss vdd d2.r_reg\[89\] _0110_ _0344_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1878_ vdd vss _0787_ _0145_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1947_ vdd vss _0793_ _0208_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_56_110 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_5_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_187 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_28_390 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1663_ vss vdd _0847_ d2.t_load\[45\] d5.fll_core.tmp\[0\] _0733_ vss vdd sky130_fd_sc_hd__mux2_1
X_1732_ vss vdd _0769_ _0017_ _0768_ vss vdd sky130_fd_sc_hd__nor2_1
X_1801_ vdd vss _0779_ _0076_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_7_261 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1594_ vss vdd _0275_ _0687_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2146_ vss vdd d2.t_load\[35\] _0162_ _0396_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2215_ vss vdd d5.fll_core.counter1.count\[3\] _0228_ _0004_ clknet_1_0__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_327 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2077_ vss vdd d2.r_reg\[72\] _0093_ _0327_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_34_360 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1028_ vss vdd _0440_ _0821_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_14_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_29_121 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_179 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_44_102 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_25_382 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_253 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2000_ vdd vss _0795_ _0250_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_35_113 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_50_149 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_16_382 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1715_ vdd vss d5.fll_core.counter1.count\[7\] d5.fll_core.counter1.count\[8\] _0760_
+ _0757_ vss vdd sky130_fd_sc_hd__a21oi_1
X_1646_ vss vdd _0706_ d2.r_reg\[3\] _0722_ _0723_ vss vdd sky130_fd_sc_hd__mux2_1
X_1577_ vss vdd _0662_ d2.r_reg\[25\] _0675_ _0676_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_58_216 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_66_293 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2129_ vss vdd d2.t_load\[18\] _0145_ _0379_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XPHY_69 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_58 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_47 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_14 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_25 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_36 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_22_341 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_66_10 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_2_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_9_323 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1500_ vss vdd _0618_ d2.r_reg\[49\] _0622_ _0623_ vss vdd sky130_fd_sc_hd__mux2_1
X_1293_ vss vdd _0463_ _0472_ _0464_ _0471_ d2.t_load\[15\] d2.t_load\[14\] vss vdd
+ sky130_fd_sc_hd__o221a_1
X_1431_ vss vdd _0326_ _0575_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1362_ vss vdd _0904_ d2.r_reg\[92\] _0527_ _0528_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_63_274 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_48_271 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_23_105 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_23_149 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1629_ vss vdd _0264_ _0711_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_11_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_46_208 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_52_78 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_45_230 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_60_277 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1980_ vdd vss _0800_ _0231_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_13_160 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_13_193 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_5_381 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1345_ vss vdd _0958_ _0516_ _0515_ vss vdd sky130_fd_sc_hd__nor2_1
X_1276_ vdd vss _0988_ d5.fll_core.counter2.count\[7\] d2.t_load\[2\] _0986_ _0985_
+ _0987_ vss vdd sky130_fd_sc_hd__a221o_1
X_1414_ vss vdd _0331_ _0563_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_51_233 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_22_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_333 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_59_300 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_0_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1130_ vss vdd _0392_ _0875_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_33_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1061_ vss vdd _0836_ d2.r_reg\[63\] d2.t_load\[63\] _0839_ vss vdd sky130_fd_sc_hd__mux2_1
X_1894_ vdd vss _0788_ _0160_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_33_299 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1963_ vdd vss _0795_ _0222_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_56_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1328_ vss vdd _0503_ d5.fll_core.tmp\[4\] _0502_ _0947_ vss vdd sky130_fd_sc_hd__a21bo_1
X_1259_ vdd vss d2.t_load\[8\] _0972_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_17_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_62_317 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2231_ vss vdd d5.fll_core.counter2.count\[9\] _0244_ _0020_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_2_181 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1113_ vss vdd _0400_ _0866_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_53_328 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_38_347 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_38_314 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2162_ vss vdd d2.t_load\[51\] _0178_ _0412_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2093_ vss vdd d2.r_reg\[88\] _0109_ _0343_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1044_ vss vdd _0825_ d2.r_reg\[71\] net22 _0830_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_17_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_61_383 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_21_225 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1877_ vdd vss _0787_ _0144_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1946_ vdd vss _0793_ _0207_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_56_133 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_62_158 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_62_125 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1800_ vdd vss _0779_ _0075_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1662_ vss vdd net7 _0732_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1731_ vss vdd _0766_ _0769_ d5.fll_core.counter2.count\[6\] vss vdd sky130_fd_sc_hd__nor2_1
X_2214_ vss vdd d5.fll_core.counter1.count\[2\] _0227_ _0003_ clknet_1_0__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1593_ vss vdd _0684_ d2.r_reg\[20\] _0686_ _0687_ vss vdd sky130_fd_sc_hd__mux2_1
X_2145_ vss vdd d2.t_load\[34\] _0161_ _0395_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_38_122 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1027_ vss vdd _0814_ d2.r_reg\[79\] net30 _0821_ vss vdd sky130_fd_sc_hd__mux2_1
X_2076_ vss vdd d2.r_reg\[71\] _0092_ _0326_ clknet_4_0_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1929_ vdd vss _0792_ _0191_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_30_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_39_57 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_17_306 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_44_136 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_265 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_35_169 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_43_191 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1714_ vss vdd _0759_ d5.fll_core.counter1.count\[7\] d5.fll_core.counter1.count\[8\]
+ _0757_ vss vdd sky130_fd_sc_hd__and3_1
X_1576_ vss vdd _0674_ d2.t_load\[25\] d2.r_reg\[26\] _0675_ vss vdd sky130_fd_sc_hd__mux2_1
X_1645_ vss vdd _0519_ d2.t_load\[3\] d2.r_reg\[4\] _0722_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_66_272 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_2128_ vss vdd d2.t_load\[17\] _0144_ _0378_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XPHY_59 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_2059_ vss vdd d2.r_reg\[54\] _0075_ _0309_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_25_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XPHY_48 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_15 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_26 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_37 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_66_22 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
Xclkbuf_1_1__f_ref_in vss vdd clknet_1_1__leaf_ref_in clknet_0_ref_in vss vdd sky130_fd_sc_hd__clkbuf_16
XFILLER_17_169 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_32_117 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1430_ vss vdd _0574_ d2.r_reg\[71\] _0573_ _0575_ vss vdd sky130_fd_sc_hd__mux2_1
X_1292_ vdd vss _0471_ _0465_ d2.t_load\[14\] d2.t_load\[13\] _0464_ _0470_ vss vdd
+ sky130_fd_sc_hd__a221o_1
X_1361_ vss vdd _0520_ net43 d2.r_reg\[93\] _0527_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_63_286 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_23_139 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_23_128 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_11_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1559_ vss vdd _0286_ _0663_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1628_ vss vdd _0706_ d2.r_reg\[9\] _0710_ _0711_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_54_253 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_14_117 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_10_345 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1413_ vss vdd _0552_ d2.r_reg\[76\] _0562_ _0563_ vss vdd sky130_fd_sc_hd__mux2_1
X_1344_ vss vdd _0946_ _0515_ _0957_ vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_3_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1275_ vdd vss d5.fll_core.counter2.count\[6\] _0987_ d2.t_load\[6\] vss vdd sky130_fd_sc_hd__xor2_1$1
XFILLER_36_275 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_47_79 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_27_286 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_63_89 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_8_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_10_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_65_359 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1060_ vss vdd _0425_ _0838_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_33_234 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1962_ vdd vss _0795_ _0221_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_18_253 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1893_ vdd vss _0788_ _0159_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1327_ vss vdd _0502_ _0964_ _0962_ vss vdd sky130_fd_sc_hd__nand2_1$1
X_1258_ vss vdd _0970_ _0971_ _0969_ vss vdd sky130_fd_sc_hd__xnor2_1$1
XFILLER_17_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1189_ vss vdd _0904_ d2.r_reg\[3\] d2.t_load\[3\] _0907_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_15_289 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_23_81 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_38_304 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2230_ vss vdd d5.fll_core.counter2.count\[8\] _0243_ _0019_ clknet_1_0__leaf_ref_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_65_101 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1112_ vss vdd _0859_ d2.r_reg\[39\] d2.t_load\[39\] _0866_ vss vdd sky130_fd_sc_hd__mux2_1
X_2161_ vss vdd d2.t_load\[50\] _0177_ _0411_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_0_85 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_0_96 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2092_ vss vdd d2.r_reg\[87\] _0108_ _0342_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1043_ vss vdd _0433_ _0829_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1945_ vdd vss _0793_ _0206_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_21_237 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1876_ vdd vss _0787_ _0143_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_56_156 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_56_123 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_56_101 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_28_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1592_ vss vdd _0674_ d2.t_load\[20\] d2.r_reg\[21\] _0686_ vss vdd sky130_fd_sc_hd__mux2_1
X_1661_ vss vdd d2.t_load\[33\] d2.t_load\[32\] d5.fll_core.corner_tmp\[2\] _0732_
+ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_50_90 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1730_ vdd vss _0768_ _0766_ d5.fll_core.counter2.count\[6\] vss vdd sky130_fd_sc_hd__and2_1$1
XFILLER_11_281 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2144_ vss vdd d2.t_load\[33\] _0160_ _0394_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_2
X_2213_ vss vdd d5.fll_core.counter1.count\[1\] _0226_ _0002_ clknet_1_0__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_2
XFILLER_38_178 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_26_318 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1026_ vss vdd _0441_ _0820_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2075_ vss vdd d2.r_reg\[70\] _0091_ _0325_ clknet_4_0_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1928_ vdd vss _0792_ _0772_ vss vdd sky130_fd_sc_hd__buf_4$1
X_1859_ vdd vss _0785_ _0128_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_29_145 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_52_181 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_40_376 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_4_277 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_50_129 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_31_310 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1713_ vss vdd _0757_ _0008_ _0473_ vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1575_ vss vdd _0674_ net2 vss vdd sky130_fd_sc_hd__clkbuf_4$1
X_1644_ vss vdd _0259_ _0721_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2127_ vss vdd d2.t_load\[16\] _0143_ _0377_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_137 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_34_181 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_2058_ vss vdd d2.r_reg\[53\] _0074_ _0308_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_159 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_25_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XPHY_49 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_16 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1009_ vss vdd _0449_ _0811_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XPHY_27 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_38 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_22_376 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_22_365 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_1_225 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_17_126 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_13_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1360_ vss vdd _0348_ _0526_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1291_ vss vdd _0465_ _0470_ _0466_ _0469_ d2.t_load\[13\] d2.t_load\[12\] vss vdd
+ sky130_fd_sc_hd__o221a_1
XFILLER_63_298 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_23_118 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1558_ vss vdd _0662_ d2.r_reg\[31\] _0661_ _0663_ vss vdd sky130_fd_sc_hd__mux2_1
X_1627_ vss vdd _0696_ d2.t_load\[9\] d2.r_reg\[10\] _0710_ vss vdd sky130_fd_sc_hd__mux2_1
X_1489_ vss vdd _0608_ d2.t_load\[52\] d2.r_reg\[53\] _0615_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_54_276 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_14_107 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_6_317 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_7_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_45_276 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_155 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1343_ vss vdd _0353_ _0514_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1412_ vss vdd _0542_ net27 d2.r_reg\[77\] _0562_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_36_243 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1274_ vdd vss d2.t_load\[7\] _0986_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_63_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_42_235 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_37_80 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1892_ vdd vss _0788_ _0158_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1961_ vss vdd _0795_ _0772_ vss vdd sky130_fd_sc_hd__clkbuf_8
X_1326_ vss vdd _0357_ _0501_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1257_ vss vdd _0946_ _0970_ d5.fll_core.tmp\[9\] vss vdd sky130_fd_sc_hd__xnor2_1$1
X_1188_ vss vdd _0365_ _0906_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_17_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_15_246 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_65_113 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_2160_ vss vdd d2.t_load\[49\] _0176_ _0410_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1111_ vss vdd _0401_ _0865_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_53_319 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2091_ vss vdd d2.r_reg\[86\] _0107_ _0341_ clknet_4_5_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_0_20 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1042_ vss vdd _0825_ d2.r_reg\[72\] net23 _0829_ vss vdd sky130_fd_sc_hd__mux2_1
Xclkbuf_4_15_0_clk_in vss vdd clknet_4_15_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
X_1875_ vdd vss _0787_ _0142_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1944_ vdd vss _0793_ _0205_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_9_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_21_205 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1309_ vss vdd _0488_ _0486_ d5.fll_core.tmp\[9\] d5.fll_core.tmp\[8\] _0487_ vss
+ vdd sky130_fd_sc_hd__and4_1
XFILLER_44_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_8_209 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_28_371 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_43_385 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_11_271 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1591_ vss vdd _0276_ _0685_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1660_ vss vdd net6 _0731_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_2212_ vss vdd d5.fll_core.counter1.count\[0\] _0225_ _0001_ clknet_1_0__leaf_vco_in
+ vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2143_ vss vdd d2.t_load\[32\] _0159_ _0393_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_38_135 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_22_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1025_ vss vdd _0814_ d2.r_reg\[80\] net31 _0820_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_14_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2074_ vss vdd d2.r_reg\[69\] _0090_ _0324_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1927_ vdd vss _0791_ _0190_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1858_ vdd vss _0785_ _0127_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1789_ vdd vss _0778_ _0065_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_39_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_69 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_29_113 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_31_333 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1712_ vss vdd _0758_ _0007_ _0757_ vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_6_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1643_ vss vdd _0706_ d2.r_reg\[4\] _0720_ _0721_ vss vdd sky130_fd_sc_hd__mux2_1
X_1574_ vss vdd _0281_ _0673_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_6_85 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_66_241 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2126_ vss vdd d2.t_load\[15\] _0142_ _0376_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2057_ vss vdd d2.r_reg\[52\] _0073_ _0307_ clknet_4_6_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_149 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XPHY_17 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XPHY_28 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_41_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_25_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1008_ vss vdd _0803_ d2.r_reg\[88\] net39 _0811_ vss vdd sky130_fd_sc_hd__mux2_1
XPHY_39 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_22_333 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_22_388 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_66_57 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_1_237 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_25_160 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_9_337 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_13_377 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1290_ vdd vss _0469_ _0467_ d2.t_load\[12\] d2.t_load\[11\] _0466_ _0468_ vss vdd
+ sky130_fd_sc_hd__a221o_1
XFILLER_48_230 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_0_281 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
Xclkbuf_4_3_0_clk_in vss vdd clknet_4_3_0_clk_in clknet_0_clk_in vss vdd sky130_fd_sc_hd__clkbuf_8
X_1626_ vss vdd _0265_ _0709_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1557_ vss vdd _0662_ _0892_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_39_241 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1488_ vss vdd _0308_ _0614_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_54_233 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_52_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2109_ vss vdd d5.fll_core.tmp\[8\] _0125_ _0359_ clknet_1_0__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_10_358 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_22_141 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_9_101 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_9_123 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1342_ vss vdd _0491_ d5.fll_core.tmp\[2\] _0513_ _0514_ vss vdd sky130_fd_sc_hd__mux2_1
X_1273_ vdd vss d5.fll_core.counter2.count\[2\] _0985_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1411_ vss vdd _0332_ _0561_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xclkbuf_0_ref_in vss vdd clknet_0_ref_in ref_in vss vdd sky130_fd_sc_hd__clkbuf_16
XFILLER_22_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1609_ vss vdd _0684_ d2.r_reg\[15\] _0697_ _0698_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_63_69 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_2_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_2_321 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_33_225 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1891_ vdd vss _0788_ _0157_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_53_91 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_33_258 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1960_ vdd vss _0794_ _0220_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_52_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1256_ vdd vss _0950_ _0948_ _0969_ _0968_ vss vdd sky130_fd_sc_hd__a21oi_1
X_1325_ vss vdd _0491_ d5.fll_core.tmp\[6\] _0500_ _0501_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_64_361 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1187_ vss vdd _0904_ d2.r_reg\[4\] d2.t_load\[4\] _0906_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_3_129 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_47_328 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_47_317 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_15_225 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_30_239 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_15_236 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1110_ vss vdd _0859_ d2.r_reg\[40\] d2.t_load\[40\] _0865_ vss vdd sky130_fd_sc_hd__mux2_1
X_2090_ vss vdd d2.r_reg\[85\] _0106_ _0340_ clknet_4_4_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_46_383 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1041_ vss vdd _0434_ _0828_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1874_ vdd vss _0787_ _0141_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1943_ vdd vss _0793_ _0204_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_44_309 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1308_ vss vdd _0487_ d5.fll_core.tmp\[5\] d5.fll_core.tmp\[7\] d5.fll_core.tmp\[6\]
+ d5.fll_core.tmp\[4\] vss vdd sky130_fd_sc_hd__and4_1
XFILLER_37_372 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1239_ vss vdd _0946_ _0952_ d5.fll_core.tmp\[7\] vss vdd sky130_fd_sc_hd__xnor2_1$1
XFILLER_29_306 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_7_210 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1590_ vss vdd _0684_ d2.r_reg\[21\] _0683_ _0685_ vss vdd sky130_fd_sc_hd__mux2_1
X_2142_ vss vdd d2.t_load\[31\] _0158_ _0392_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2211_ vdd vss d5.fll_core.corner_tmp\[2\] clknet_1_1__leaf_ref_in _0459_ vss vdd
+ sky130_fd_sc_hd__dfxtp_1
X_2073_ vss vdd d2.r_reg\[68\] _0089_ _0323_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1024_ vss vdd _0442_ _0819_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_15_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_46_180 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1788_ vdd vss _0778_ _0064_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1926_ vdd vss _0791_ _0189_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1857_ vdd vss _0785_ _0126_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_30_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_39_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_37_191 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_29_158 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_25_375 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_25_331 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_345 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_40_334 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_4_213 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_62 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_28_180 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1711_ vss vdd _0755_ _0758_ d5.fll_core.counter1.count\[6\] vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_6_20 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_6_53 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1642_ vss vdd _0519_ d2.t_load\[4\] d2.r_reg\[5\] _0720_ vss vdd sky130_fd_sc_hd__mux2_1
X_1573_ vss vdd _0662_ d2.r_reg\[26\] _0672_ _0673_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_58_209 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_6_97 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2125_ vss vdd d2.t_load\[14\] _0141_ _0375_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2056_ vss vdd d2.r_reg\[51\] _0072_ _0306_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_117 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XPHY_18 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1007_ vss vdd _0450_ _0810_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XPHY_29 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_22_301 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1909_ vdd vss _0790_ _0173_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_41_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_1_205 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_49_209 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_15_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_197 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_63_212 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_48_264 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_0_293 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1556_ vss vdd _0652_ d2.t_load\[31\] d2.r_reg\[32\] _0661_ vss vdd sky130_fd_sc_hd__mux2_1
X_1625_ vss vdd _0706_ d2.r_reg\[10\] _0708_ _0709_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_8_360 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1487_ vss vdd _0596_ d2.r_reg\[53\] _0613_ _0614_ vss vdd sky130_fd_sc_hd__mux2_1
X_2039_ vss vdd d2.r_reg\[34\] _0055_ _0289_ clknet_4_11_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2108_ vss vdd d5.fll_core.tmp\[7\] _0124_ _0358_ clknet_1_0__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_22_153 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_22_197 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_45_289 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_9_113 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1410_ vss vdd _0552_ d2.r_reg\[77\] _0560_ _0561_ vss vdd sky130_fd_sc_hd__mux2_1
X_1341_ vdd vss _0960_ _0513_ _0955_ vss vdd sky130_fd_sc_hd__xor2_1$1
X_1272_ vdd vss d2.t_load\[4\] _0984_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_51_215 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1539_ vss vdd _0292_ _0649_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_59_326 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1608_ vss vdd _0696_ d2.t_load\[15\] d2.r_reg\[16\] _0697_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_63_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_59_359 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_10_178 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_12_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_12_85 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_2_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_2_333 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_33_215 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1890_ vdd vss _0788_ _0156_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_45_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_49_370 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1255_ vss vdd _0968_ _0965_ _0947_ _0967_ _0953_ _0962_ vss vdd sky130_fd_sc_hd__a32o_1
X_1324_ vdd vss _0495_ _0500_ _0951_ vss vdd sky130_fd_sc_hd__xor2_1$1
X_1186_ vss vdd _0366_ _0905_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_58_15 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_47_307 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_30_229 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_23_292 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_174 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_141 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_65_148 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_48_81 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1040_ vss vdd _0825_ d2.r_reg\[73\] net24 _0828_ vss vdd sky130_fd_sc_hd__mux2_1
X_1942_ vdd vss _0793_ _0203_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1873_ vdd vss _0787_ _0780_ vss vdd sky130_fd_sc_hd__buf_4$1
XFILLER_28_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1307_ vss vdd _0486_ d5.fll_core.tmp\[1\] d5.fll_core.tmp\[2\] d5.fll_core.tmp\[0\]
+ vss vdd sky130_fd_sc_hd__and3_1
X_1169_ vss vdd _0374_ _0896_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1238_ vss vdd _0946_ _0951_ d5.fll_core.tmp\[6\] vss vdd sky130_fd_sc_hd__xnor2_1$1
XFILLER_52_365 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_7_299 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2210_ vdd vss d5.fll_core.corner_tmp\[1\] clknet_1_1__leaf_ref_in _0458_ vss vdd
+ sky130_fd_sc_hd__dfxtp_1
X_2141_ vss vdd d2.t_load\[30\] _0157_ _0391_ clknet_4_15_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_53_118 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2072_ vss vdd d2.r_reg\[67\] _0088_ _0322_ clknet_4_3_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1023_ vss vdd _0814_ d2.r_reg\[81\] net32 _0819_ vss vdd sky130_fd_sc_hd__mux2_1
X_1925_ vdd vss _0791_ _0188_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_34_376 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1787_ vdd vss _0778_ _0063_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1856_ vdd vss _0785_ _0125_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_39_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_96 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_16_332 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1572_ vss vdd _0652_ d2.t_load\[26\] d2.r_reg\[27\] _0672_ vss vdd sky130_fd_sc_hd__mux2_1
X_1710_ vdd vss _0757_ _0755_ d5.fll_core.counter1.count\[6\] vss vdd sky130_fd_sc_hd__and2_1$1
XFILLER_6_65 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1641_ vss vdd _0260_ _0719_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_66_221 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_2124_ vss vdd d2.t_load\[13\] _0140_ _0374_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_66_265 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2055_ vss vdd d2.r_reg\[50\] _0071_ _0305_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_26_107 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XPHY_19 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1006_ vss vdd _0803_ d2.r_reg\[89\] net40 _0810_ vss vdd sky130_fd_sc_hd__mux2_1
X_1908_ vdd vss _0790_ _0172_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1839_ vdd vss _0783_ _0110_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_57_254 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_154 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xoutput5 vss vdd corner[0] net5 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_31_95 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_31_51 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xoutput40 vss vdd vbias3[4] net40 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_56_81 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1555_ vss vdd _0287_ _0660_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1624_ vss vdd _0696_ d2.t_load\[10\] d2.r_reg\[11\] _0708_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_54_202 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_36_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_2107_ vss vdd d5.fll_core.tmp\[6\] _0123_ _0357_ clknet_1_0__leaf_ref_in vss vdd
+ sky130_fd_sc_hd__dfrtp_2
X_1486_ vss vdd _0608_ d2.t_load\[53\] d2.r_reg\[54\] _0613_ vss vdd sky130_fd_sc_hd__mux2_1
X_2038_ vss vdd d2.r_reg\[33\] _0054_ _0288_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
XFILLER_54_246 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_10_305 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_22_165 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_6_309 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_9_169 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_54_8 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1340_ vss vdd _0354_ _0512_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1271_ vss vdd _0983_ d5.fll_core.counter2.count\[8\] _0976_ _0972_ _0982_ vss vdd
+ sky130_fd_sc_hd__a211o_1
X_1538_ vss vdd _0640_ d2.r_reg\[37\] _0648_ _0649_ vss vdd sky130_fd_sc_hd__mux2_1
X_1469_ vss vdd _0314_ _0601_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1607_ vss vdd _0696_ net2 vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_63_27 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_10_146 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_10_168 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_5_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_2_345 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_2_389 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_279 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_41_293 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_41_271 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_38_3 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1323_ vss vdd _0358_ _0499_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_49_382 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1254_ vdd vss d5.fll_core.tmp\[7\] _0967_ d5.fll_core.tmp\[6\] _0966_ vss vdd sky130_fd_sc_hd__or3_1
X_1185_ vss vdd _0904_ d2.r_reg\[5\] d2.t_load\[5\] _0905_ vss vdd sky130_fd_sc_hd__mux2_1
XFILLER_59_124 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_55_363 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_55_330 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_30_219 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_2_197 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_0_67 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_61_333 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
X_1872_ vdd vss _0786_ _0140_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1941_ vdd vss _0793_ _0202_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1306_ vdd vss _0961_ _0956_ _0485_ _0967_ _0484_ vss vdd sky130_fd_sc_hd__or4_1
XFILLER_52_377 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_52_344 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
X_1099_ vss vdd _0859_ _0802_ vss vdd sky130_fd_sc_hd__clkbuf_4$1
XFILLER_44_29 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1168_ vss vdd _0893_ d2.r_reg\[13\] d2.t_load\[13\] _0896_ vss vdd sky130_fd_sc_hd__mux2_1
X_1237_ vss vdd _0949_ _0950_ _0948_ vss vdd sky130_fd_sc_hd__nor2_1
XFILLER_20_241 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_20_274 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_47_138 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_41 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_43_322 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_18_96 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_11_296 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_2140_ vss vdd d2.t_load\[29\] _0156_ _0390_ clknet_4_14_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2071_ vss vdd d2.r_reg\[66\] _0087_ _0321_ clknet_4_2_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1022_ vss vdd _0443_ _0818_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1924_ vdd vss _0791_ _0187_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1855_ vdd vss _0785_ _0124_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_34_388 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1786_ vdd vss _0778_ _0062_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_55_39 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_52_141 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_25_344 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_20_20 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_20_53 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_61_93 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_31_325 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_31_303 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
X_1571_ vss vdd _0282_ _0671_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_3_281 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_6_77 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
X_1640_ vss vdd _0706_ d2.r_reg\[5\] _0718_ _0719_ vss vdd sky130_fd_sc_hd__mux2_1
X_2123_ vss vdd d2.t_load\[12\] _0139_ _0373_ clknet_4_13_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_2054_ vss vdd d2.r_reg\[49\] _0070_ _0304_ clknet_4_12_0_clk_in vss vdd sky130_fd_sc_hd__dfrtp_1$1
X_1005_ vss vdd _0451_ _0809_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_19_182 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1907_ vdd vss _0790_ _0171_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1838_ vdd vss _0783_ _0109_ vss vdd sky130_fd_sc_hd__inv_2$1
X_1769_ vdd vss _0776_ _0047_ vss vdd sky130_fd_sc_hd__inv_2$1
XFILLER_57_211 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
XFILLER_1_218 vdd vss vss vdd sky130_fd_sc_hd__decap_6$1
XFILLER_57_299 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_40_188 vdd vss vss vdd sky130_fd_sc_hd__decap_8$1
XFILLER_25_196 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_25_152 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
XFILLER_15_75 vss vdd vss vdd sky130_fd_sc_hd__decap_4$1
Xoutput6 vss vdd corner[1] net6 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput41 vss vdd vbias3[5] net41 vss vdd sky130_fd_sc_hd__clkbuf_1$1
Xoutput30 vss vdd vbias2[2] net30 vss vdd sky130_fd_sc_hd__clkbuf_1$1
XFILLER_63_225 vdd vss vss vdd sky130_fd_sc_hd__decap_3$1
XFILLER_16_141 vss vdd vss vdd sky130_ef_sc_hd__decap_12$1
X_1554_ vss vdd _0640_ d2.r_reg\[32\] _0659_ _0660_ vss vdd sky130_fd_sc_hd__mux2_1
X_1623_ vss vdd _0266_ _0707_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
X_1485_ vss vdd _0309_ _0612_ vss vdd sky130_fd_sc_hd__clkbuf_1$1
.ends

.subckt o_n_3 a_159_n70# a_n707_n244# a_351_n70# a_n33_n70# a_n225_n70# a_n465_92#
+ a_n417_n70#
X0 a_n707_n244# a_n465_92# a_n33_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n33_n70# a_n465_92# a_n707_n244# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_159_n70# a_n465_92# a_n707_n244# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n707_n244# a_n465_92# a_159_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_351_n70# a_n465_92# a_n707_n244# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n707_n244# a_n465_92# a_351_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X6 a_n707_n244# a_n707_n244# a_n707_n244# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 a_n707_n244# a_n465_92# a_n417_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X8 a_n707_n244# a_n707_n244# a_n707_n244# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X9 a_n417_n70# a_n465_92# a_n707_n244# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X10 a_n225_n70# a_n465_92# a_n707_n244# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X11 a_n707_n244# a_n465_92# a_n225_n70# a_n707_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt o_p_1 w_n1319_n289# a_n1041_n167# a_n993_n70#
X0 a_n1041_n167# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 w_n1319_n289# a_n1041_n167# a_n1041_n167# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 w_n1319_n289# w_n1319_n289# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X6 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X8 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X9 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X10 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X11 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X12 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X13 w_n1319_n289# w_n1319_n289# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X14 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X15 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X16 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X17 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X18 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X19 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X20 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X21 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X22 a_n993_n70# a_n1041_n167# w_n1319_n289# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X23 w_n1319_n289# a_n1041_n167# a_n993_n70# w_n1319_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt o_n_2 a_n221_n70# a_n33_n70# a_n323_n244# a_n81_n158#
X0 a_n221_n70# a_n81_n158# a_n33_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n33_n70# a_n81_n158# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n221_n70# a_n221_n70# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n221_n70# a_n221_n70# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt ota_half sky130_fd_pr__pfet_01v8_BDSGKN_0/a_n1041_n167# sky130_fd_pr__nfet_01v8_CCWHWC_0/a_n417_n70#
+ sky130_fd_pr__nfet_01v8_CCWHWC_0/a_159_n70# sky130_fd_pr__nfet_01v8_2AA63J_0/a_n221_n70#
+ sky130_fd_pr__nfet_01v8_2AA63J_0/a_n33_n70# sky130_fd_pr__nfet_01v8_CCWHWC_0/a_351_n70#
+ sky130_fd_pr__nfet_01v8_CCWHWC_0/a_n33_n70# sky130_fd_pr__nfet_01v8_CCWHWC_0/a_n465_92#
+ sky130_fd_pr__nfet_01v8_2AA63J_0/a_n81_n158# sky130_fd_pr__nfet_01v8_CCWHWC_0/a_n225_n70#
+ sky130_fd_pr__pfet_01v8_BDSGKN_0/w_n1319_n289# VSUBS sky130_fd_pr__pfet_01v8_BDSGKN_0/a_n993_n70#
Xsky130_fd_pr__nfet_01v8_CCWHWC_0 sky130_fd_pr__nfet_01v8_CCWHWC_0/a_159_n70# VSUBS
+ sky130_fd_pr__nfet_01v8_CCWHWC_0/a_351_n70# sky130_fd_pr__nfet_01v8_CCWHWC_0/a_n33_n70#
+ sky130_fd_pr__nfet_01v8_CCWHWC_0/a_n225_n70# sky130_fd_pr__nfet_01v8_CCWHWC_0/a_n465_92#
+ sky130_fd_pr__nfet_01v8_CCWHWC_0/a_n417_n70# o_n_3
Xsky130_fd_pr__pfet_01v8_BDSGKN_0 sky130_fd_pr__pfet_01v8_BDSGKN_0/w_n1319_n289# sky130_fd_pr__pfet_01v8_BDSGKN_0/a_n1041_n167#
+ sky130_fd_pr__pfet_01v8_BDSGKN_0/a_n993_n70# o_p_1
Xsky130_fd_pr__nfet_01v8_2AA63J_0 sky130_fd_pr__nfet_01v8_2AA63J_0/a_n221_n70# sky130_fd_pr__nfet_01v8_2AA63J_0/a_n33_n70#
+ VSUBS sky130_fd_pr__nfet_01v8_2AA63J_0/a_n81_n158# o_n_2
.ends

.subckt ota_bias a_n273_92# a_n515_n244# a_n225_n70#
X0 a_n515_n244# a_n273_92# a_n225_n70# a_n515_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n225_n70# a_n273_92# a_n515_n244# a_n515_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n225_n70# a_n273_92# a_n515_n244# a_n515_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n515_n244# a_n273_92# a_n225_n70# a_n515_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n515_n244# a_n515_n244# a_n515_n244# a_n515_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n515_n244# a_n515_n244# a_n515_n244# a_n515_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X6 a_n225_n70# a_n273_92# a_n515_n244# a_n515_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 a_n515_n244# a_n273_92# a_n225_n70# a_n515_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt ota_2 in_p in_n vbias vdd out net1 vss
Xota_half_0 m1_2226_350# m1_609_381# m1_609_381# net1 m1_2226_350# m1_609_381# m1_609_381#
+ m1_609_381# in_n m1_609_381# vdd vss m1_609_381# ota_half
Xota_half_1 m1_3004_350# out out net1 m1_3004_350# out out m1_609_381# in_p out vdd
+ vss out ota_half
Xota_bias_0 vbias vss net1 ota_bias
.ends

.subckt diff_p w_n455_n289# a_n317_n70# a_n129_n70# a_n177_n167#
X0 a_n317_n70# a_n177_n167# a_n129_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n317_n70# a_n177_n167# a_n129_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n317_n70# a_n317_n70# a_n317_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n317_n70# a_n317_n70# a_n317_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n129_n70# a_n177_n167# a_n317_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n129_n70# a_n177_n167# a_n317_n70# w_n455_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt diff_n a_n221_n70# a_n81_92# a_n33_n70# a_n323_n244#
X0 a_n221_n70# a_n81_92# a_n33_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n33_n70# a_n81_92# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n221_n70# a_n221_n70# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n221_n70# a_n221_n70# a_n221_n70# a_n323_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt differential clk_in nclk clk vdd vss
Xdiff_p_0 vdd m2_772_1987# inv_simple1_3/in clk_in diff_p
Xdiff_n_0 m2_1060_1348# clk_in inv_simple1_3/in vss diff_n
Xsky130_fd_pr__pfet_01v8_X6FFBL_0 vdd m2_772_1987# vdd vss diff_p
Xinv_simple1_0 clk_in inv_simple1_1/in vdd vss inv_simple1
Xinv_simple1_1 inv_simple1_1/in inv_simple1_2/in vdd vss inv_simple1
Xinv_simple1_3 inv_simple1_3/in clk vdd vss inv_simple1
Xinv_simple1_2 inv_simple1_2/in nclk vdd vss inv_simple1
Xsky130_fd_pr__nfet_01v8_2AA63J_0 m2_1060_1348# vdd vss vss diff_n
.ends

.subckt cap50f c1_n550_n500# m3_n650_n600#
X0 c1_n550_n500# m3_n650_n600# sky130_fd_pr__cap_mim_m3_1 l=5e+06u w=5e+06u
.ends

.subckt sspd ref_in vco_in vbias v_out vdd vss
Xota_2_0 ota_2_0/in_p ota_2_0/out vbias vdd ota_2_0/out ota_2_0/net1 vss ota_2
Xinv_buffer2_0 ref_in inv_buffer2_0/out1 vdd vss inv_buffer2
Xdifferential_0 inv_buffer2_0/out1 tgate_1_0/sw tgate_1_1/sw vdd vss differential
Xtgate_1_1 tgate_1_1/sw v_out vdd vss ota_2_0/out tgate_1
Xtgate_1_0 tgate_1_0/sw ota_2_0/in_p vdd vss vco_in tgate_1
Xcap50f_0 ota_2_0/in_p vss cap50f
.ends

.subckt cap_200p m3_n3186_n3040# c1_n3146_n3000#
X0 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X1 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X2 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X3 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X4 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X5 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X6 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X7 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X8 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X9 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X10 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X11 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X12 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X13 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X14 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X15 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X16 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X17 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X18 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X19 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X20 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X21 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X22 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X23 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X24 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X25 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X26 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X27 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X28 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X29 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X30 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X31 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X32 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X33 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X34 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X35 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X36 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X37 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X38 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X39 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X40 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X41 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X42 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X43 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X44 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X45 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X46 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X47 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X48 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X49 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X50 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X51 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X52 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X53 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X54 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X55 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X56 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X57 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X58 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X59 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X60 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X61 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X62 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X63 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X64 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X65 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X66 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X67 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X68 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X69 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X70 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X71 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X72 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X73 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X74 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X75 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X76 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X77 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X78 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X79 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X80 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X81 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X82 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X83 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X84 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X85 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X86 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X87 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X88 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X89 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X90 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X91 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X92 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X93 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X94 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X95 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X96 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X97 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X98 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X99 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X100 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X101 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X102 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X103 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X104 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X105 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X106 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X107 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X108 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
X109 c1_n3146_n3000# m3_n3186_n3040# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=3e+07u
.ends

.subckt r_8k a_942_1771# vss a_n1512_1771#
X0 a_n1512_n2203# a_n1512_1771# vss sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X1 a_124_n2203# a_n694_1771# vss sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X2 a_n1512_n2203# a_n694_1771# vss sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X3 vss vss vss sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X4 a_124_n2203# a_942_1771# vss sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
X5 vss vss vss sky130_fd_pr__res_high_po w=2.85e+06u l=1.771e+07u
.ends

.subckt voltage_control vcoarse vfine vdd vout lock vss
Xcap_200p_0 vout vss cap_200p
Xr_8k_0 vout vss vcoarse r_8k
Xinv_simple1_0 lock tgate_1_0/sw vdd vss inv_simple1
Xtgate_1_0 tgate_1_0/sw vcoarse vdd vss vfine tgate_1
.ends

.subckt stf_ctrl vctrl swff swtt swss b0 b1 b2 vdd vss
Xtgate_1_1 vctrl swtt vdd vss b1 tgate_1
Xtgate_1_0 vctrl swss vdd vss b2 tgate_1
Xtgate_1_2 vctrl swff vdd vss b0 tgate_1
.ends

.subckt sky130_fd_sc_hd__dfxbp_1 VGND VPWR Q_N D CLK Q VNB VPB
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X4 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X9 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VGND a_1059_315# a_1490_369# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=750000u l=150000u
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X17 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X19 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=360000u l=150000u
X21 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
X22 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 Q_N a_1490_369# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X25 Q_N a_1490_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X27 VPWR a_1059_315# a_1490_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=640000u l=150000u
.ends

.subckt sky130_fd_sc_hd__nand2_1 VGND VPWR Y B A VNB VPB
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 Y A a_113_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 a_113_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt d_ff_15 f_15 vss vdd f_in
Xsky130_fd_sc_hd__dfxbp_1_0 vss vdd sky130_fd_sc_hd__dfxbp_1_0/Q_N sky130_fd_sc_hd__nand2_1_0/Y
+ f_in sky130_fd_sc_hd__dfxbp_1_1/D vss vdd sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__dfxbp_1_1 vss vdd sky130_fd_sc_hd__dfxbp_1_1/Q_N sky130_fd_sc_hd__dfxbp_1_1/D
+ f_in sky130_fd_sc_hd__nand2_1_0/B vss vdd sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__dfxbp_1_2 vss vdd sky130_fd_sc_hd__dfxbp_1_2/Q_N sky130_fd_sc_hd__nand2_1_0/B
+ f_in sky130_fd_sc_hd__nand2_1_0/A vss vdd sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__dfxbp_1_3 vss vdd sky130_fd_sc_hd__dfxbp_1_3/Q_N sky130_fd_sc_hd__nand2_1_1/Y
+ sky130_fd_sc_hd__dfxbp_1_1/D sky130_fd_sc_hd__nand2_1_1/B vss vdd sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__dfxbp_1_4 vss vdd f_15 sky130_fd_sc_hd__nand2_1_1/B sky130_fd_sc_hd__dfxbp_1_1/D
+ sky130_fd_sc_hd__nand2_1_1/A vss vdd sky130_fd_sc_hd__dfxbp_1
Xsky130_fd_sc_hd__nand2_1_0 vss vdd sky130_fd_sc_hd__nand2_1_0/Y sky130_fd_sc_hd__nand2_1_0/B
+ sky130_fd_sc_hd__nand2_1_0/A vss vdd sky130_fd_sc_hd__nand2_1
Xsky130_fd_sc_hd__nand2_1_1 vss vdd sky130_fd_sc_hd__nand2_1_1/Y sky130_fd_sc_hd__nand2_1_1/B
+ sky130_fd_sc_hd__nand2_1_1/A vss vdd sky130_fd_sc_hd__nand2_1
.ends

.subckt n_cell_1 a_n419_n244# a_n177_n158# a_63_n70# a_n317_n70# a_n129_n70# a_33_n158#
X0 a_63_n70# a_33_n158# a_n317_n70# a_n419_n244# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n317_n70# a_n177_n158# a_n129_n70# a_n419_n244# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n317_n70# a_n317_n70# a_n317_n70# a_n419_n244# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n317_n70# a_33_n158# a_63_n70# a_n419_n244# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n317_n70# a_n317_n70# a_n317_n70# a_n419_n244# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 a_n129_n70# a_n177_n158# a_n317_n70# a_n419_n244# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt p_cell_3 a_n321_n70# a_207_n167# a_n81_101# w_n551_n289# a_n273_101#
X0 w_n551_n289# a_n81_101# a_n321_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 w_n551_n289# w_n551_n289# a_n81_101# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 w_n551_n289# a_n81_101# a_n81_101# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 a_n81_101# a_207_n167# w_n551_n289# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 a_n321_n70# w_n551_n289# w_n551_n289# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 w_n551_n289# a_n273_101# a_n321_n70# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X6 a_n321_n70# a_n321_n70# w_n551_n289# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 a_n81_101# a_n321_n70# w_n551_n289# w_n551_n289# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt current_tails_1 swss swtt swff in vss
X0 vss swss in vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 in swss vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 in swtt vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 vss swtt in vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X4 in swtt vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X5 vss swff in vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X6 vss vss vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X7 vss swss in vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X8 vss vss vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X9 in swss vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X10 in swss vss vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X11 vss swss in vss sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt n_cell_3 a_n32_92# a_16_n70# a_n274_n244#
X0 a_16_n70# a_n32_92# a_n274_n244# a_n274_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n274_n244# a_n274_n244# a_n274_n244# a_n274_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 a_n274_n244# a_n274_n244# a_16_n70# a_n274_n244# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt sky130_fd_pr__pfet_01v8_X679XQ a_n32_n70# a_n80_101# w_n358_n288#
X0 w_n358_n288# a_n80_101# a_n32_n70# w_n358_n288# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X1 a_n32_n70# a_n80_101# w_n358_n288# w_n358_n288# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X2 w_n358_n288# w_n358_n288# w_n358_n288# w_n358_n288# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
X3 w_n358_n288# w_n358_n288# w_n358_n288# w_n358_n288# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=700000u l=150000u
.ends

.subckt delay_cell_4 din1 din2 dout1 dout2 vb b1 b0 b2 inv1 inv2 current_tails_1_0/in
+ vdd vss
Xsky130_fd_pr__nfet_01v8_lvt_GVQ53W_0 vss din1 dout2 current_tails_1_0/in dout1 din2
+ n_cell_1
Xsky130_fd_pr__pfet_01v8_X6PFBL_0 dout1 vb dout2 vdd vb p_cell_3
Xcurrent_tails_1_0 b2 b1 b0 current_tails_1_0/in vss current_tails_1
Xn_cell_3_0 vss n_cell_3_0/a_16_n70# vss n_cell_3
Xsky130_fd_pr__nfet_01v8_5ZA63U_0 dout1 inv1 vss n_cell_3
Xsky130_fd_pr__nfet_01v8_5ZA63U_1 dout2 inv2 vss n_cell_3
Xsky130_fd_pr__pfet_01v8_X679XQ_0 inv1 dout1 vdd sky130_fd_pr__pfet_01v8_X679XQ
Xsky130_fd_pr__pfet_01v8_X679XQ_1 inv2 dout2 vdd sky130_fd_pr__pfet_01v8_X679XQ
Xsky130_fd_pr__pfet_01v8_X679XQ_2 n_cell_3_0/a_16_n70# vss vdd sky130_fd_pr__pfet_01v8_X679XQ
.ends

.subckt vco_core_8 b2 b1 b0 vdelay inv1 inv2 inv3 inv4 inv5 inv6 inv7 inv8 vdd out1
+ out2 out4 out3 out7 out8 out5 out6 vss
Xdelay_cell_4_0 out8 out7 out1 out2 vdelay b1 b0 b2 inv1 inv2 delay_cell_4_0/current_tails_1_0/in
+ vdd vss delay_cell_4
Xdelay_cell_4_1 out2 out1 out3 out4 vdelay b1 b0 b2 inv4 inv3 delay_cell_4_1/current_tails_1_0/in
+ vdd vss delay_cell_4
Xdelay_cell_4_3 out6 out5 out7 out8 vdelay b1 b0 b2 inv8 inv7 delay_cell_4_3/current_tails_1_0/in
+ vdd vss delay_cell_4
Xdelay_cell_4_2 out3 out4 out5 out6 vdelay b1 b0 b2 inv5 inv6 delay_cell_4_2/current_tails_1_0/in
+ vdd vss delay_cell_4
.ends

.subckt full_vco_1 out3 out4 vbias out1 out2 b0 b1 b2 vdelay vdd vss
Xstf_ctrl_0 vbias vco_core_8_0/b0 vco_core_8_0/b1 vco_core_8_0/b2 b0 b1 b2 vdd vss
+ stf_ctrl
Xinv_buffer2_0 inv_simple1_0/out d_ff_15_0/f_in vdd vss inv_buffer2
Xinv_buffer2_1 inv_simple1_3/out d_ff_15_1/f_in vdd vss inv_buffer2
Xinv_buffer2_2 inv_simple1_6/out d_ff_15_3/f_in vdd vss inv_buffer2
Xinv_buffer2_3 inv_simple1_5/out d_ff_15_2/f_in vdd vss inv_buffer2
Xinv_simple1_0 inv_simple1_0/in inv_simple1_0/out vdd vss inv_simple1
Xd_ff_15_0 out2 vss vdd d_ff_15_0/f_in d_ff_15
Xinv_simple1_1 inv_simple1_1/in inv_simple1_1/out vdd vss inv_simple1
Xd_ff_15_1 out1 vss vdd d_ff_15_1/f_in d_ff_15
Xinv_simple1_2 inv_simple1_2/in inv_simple1_2/out vdd vss inv_simple1
Xinv_simple1_3 inv_simple1_3/in inv_simple1_3/out vdd vss inv_simple1
Xd_ff_15_2 out4 vss vdd d_ff_15_2/f_in d_ff_15
Xinv_simple1_4 inv_simple1_4/in inv_simple1_4/out vdd vss inv_simple1
Xd_ff_15_3 out3 vss vdd d_ff_15_3/f_in d_ff_15
Xvco_core_8_0 vco_core_8_0/b2 vco_core_8_0/b1 vco_core_8_0/b0 vdelay inv_simple1_3/in
+ inv_simple1_2/in inv_simple1_0/in inv_simple1_1/in inv_simple1_6/in inv_simple1_7/in
+ inv_simple1_4/in inv_simple1_5/in vdd vco_core_8_0/out1 vco_core_8_0/out2 vco_core_8_0/out4
+ vco_core_8_0/out3 vco_core_8_0/out7 vco_core_8_0/out8 vco_core_8_0/out5 vco_core_8_0/out6
+ vss vco_core_8
Xinv_simple1_5 inv_simple1_5/in inv_simple1_5/out vdd vss inv_simple1
Xinv_simple1_6 inv_simple1_6/in inv_simple1_6/out vdd vss inv_simple1
Xinv_simple1_7 inv_simple1_7/in inv_simple1_7/out vdd vss inv_simple1
.ends

.subckt full_IC_1 ref_in out vdd reset clk_in read load s_in s_out vss
Xr2r_8_0 r2r_8_0/vout r2r_8_0/b0 r2r_8_0/b1 r2r_8_0/b2 r2r_8_0/b3 r2r_8_0/b4 r2r_8_0/b5
+ r2r_8_0/b6 r2r_8_0/b7 vss r2r_8
Xr2r_8_1 sspd_0/vbias r2r_8_1/b0 r2r_8_1/b1 r2r_8_1/b2 r2r_8_1/b3 r2r_8_1/b4 r2r_8_1/b5
+ r2r_8_1/b6 r2r_8_1/b7 vss r2r_8
Xr2r_8_2 r2r_8_2/vout r2r_8_2/b0 r2r_8_2/b1 r2r_8_2/b2 r2r_8_2/b3 r2r_8_2/b4 r2r_8_2/b5
+ r2r_8_2/b6 r2r_8_2/b7 vss r2r_8
Xinv_buffer2_0 inv_buffer2_0/in1 sspd_0/ref_in vdd vss inv_buffer2
Xslopebuf_0 slopebuf_0/bit1 slopebuf_0/bit0 slopebuf_0/bit2 slopebuf_0/clk_in sspd_0/vco_in
+ vdd r2r_8_2/vout vss slopebuf
Xr2r_10_0 r2r_10_0/b0 r2r_10_0/b1 r2r_10_0/b2 r2r_10_0/b3 r2r_10_0/b4 r2r_10_0/b5
+ r2r_10_0/b6 r2r_10_0/b7 r2r_10_0/vout r2r_10_0/b8 r2r_10_0/b9 vss r2r_10
Xwrapper_0 clk_in r2r_10_0/b0 r2r_10_0/b1 r2r_10_0/b2 r2r_10_0/b3 r2r_10_0/b4 r2r_10_0/b5
+ r2r_10_0/b6 r2r_10_0/b7 load read wrapper_0/ref_in reset s_in s_out r2r_8_2/b0 r2r_8_2/b1
+ r2r_8_2/b2 r2r_8_2/b3 r2r_8_2/b4 r2r_8_2/b5 r2r_8_2/b6 r2r_8_2/b7 wrapper_0/vco_in
+ wrapper_0/_0001_ wrapper_0/_0002_ wrapper_0/_0006_ wrapper_0/_0010_ wrapper_0/_0225_
+ wrapper_0/_0226_ wrapper_0/_0227_ wrapper_0/_0229_ wrapper_0/_0230_ wrapper_0/_0463_
+ wrapper_0/_0464_ wrapper_0/_0470_ wrapper_0/_0473_ wrapper_0/_0480_ wrapper_0/_0730_
+ wrapper_0/_0732_ wrapper_0/_0751_ wrapper_0/_0752_ wrapper_0/_0753_ wrapper_0/_0754_
+ wrapper_0/_0755_ wrapper_0/_0757_ wrapper_0/_0760_ wrapper_0/_0798_ wrapper_0/_0800_
+ wrapper_0/_0912_ wrapper_0/_0913_ wrapper_0/_0914_ wrapper_0/_0915_ wrapper_0/_0918_
+ wrapper_0/_0919_ wrapper_0/_0920_ wrapper_0/_0921_ wrapper_0/_0923_ wrapper_0/_0925_
+ wrapper_0/_0930_ wrapper_0/_0931_ wrapper_0/_0932_ wrapper_0/_0936_ wrapper_0/_0938_
+ wrapper_0/_0939_ wrapper_0/_0940_ wrapper_0/_0941_ wrapper_0/_0942_ wrapper_0/_0943_
+ wrapper_0/d2.t_load\[13\] wrapper_0/d2.t_load\[25\] wrapper_0/d5.fll_core.counter1.count\[0\]
+ wrapper_0/d5.fll_core.counter1.count\[1\] wrapper_0/d5.fll_core.counter1.count\[2\]
+ wrapper_0/d5.fll_core.counter1.count\[4\] wrapper_0/d5.fll_core.counter1.count\[5\]
+ wrapper_0/d5.fll_core.counter1.count\[6\] wrapper_0/d5.fll_core.counter1.count\[7\]
+ wrapper_0/d5.fll_core.counter1.count\[8\] wrapper_0/d5.fll_core.counter_reset r2r_10_0/b9
+ wrapper_0/lock wrapper_0/net6 wrapper_0/net7 wrapper_0/_0045_ wrapper_0/_0146_ wrapper_0/_0275_
+ wrapper_0/_0276_ wrapper_0/_0787_ wrapper_0/_0788_ wrapper_0/_0277_ wrapper_0/_0278_
+ wrapper_0/_0870_ wrapper_0/_0875_ wrapper_0/_0878_ wrapper_0/_0881_ wrapper_0/_0882_
+ wrapper_0/_0883_ wrapper_0/_0884_ wrapper_0/_0885_ wrapper_0/_0886_ wrapper_0/_0888_
+ wrapper_0/_0282_ wrapper_0/_0381_ wrapper_0/_0383_ wrapper_0/_0384_ wrapper_0/_0388_
+ wrapper_0/_0389_ wrapper_0/_0147_ wrapper_0/_0148_ wrapper_0/_0465_ wrapper_0/_0467_
+ wrapper_0/_0927_ wrapper_0/_0468_ wrapper_0/_0469_ wrapper_0/_0149_ wrapper_0/_0934_
+ wrapper_0/_0150_ wrapper_0/_0937_ wrapper_0/_0151_ wrapper_0/_0652_ wrapper_0/_0671_
+ wrapper_0/_0672_ wrapper_0/_0673_ wrapper_0/_0674_ wrapper_0/clknet_4_15_0_clk_in
+ wrapper_0/d2.r_reg\[21\] wrapper_0/d2.r_reg\[22\] wrapper_0/d2.r_reg\[24\] wrapper_0/d2.r_reg\[25\]
+ wrapper_0/d2.r_reg\[27\] wrapper_0/d2.r_reg\[28\] wrapper_0/d2.r_reg\[31\] wrapper_0/_0675_
+ wrapper_0/d2.t_load\[19\] wrapper_0/d2.t_load\[20\] wrapper_0/d2.t_load\[21\] wrapper_0/d2.t_load\[23\]
+ wrapper_0/d2.t_load\[24\] wrapper_0/_0677_ wrapper_0/d2.t_load\[27\] wrapper_0/d2.t_load\[28\]
+ wrapper_0/d2.t_load\[30\] wrapper_0/d2.t_load\[31\] wrapper_0/_0678_ wrapper_0/_0679_
+ wrapper_0/_0681_ wrapper_0/_0683_ wrapper_0/_0684_ wrapper_0/_0685_ wrapper_0/_0686_
+ wrapper_0/_0689_ wrapper_0/_0154_ r2r_10_0/b8 wrapper_0/_0158_ wrapper_0/_0042_
+ wrapper_0/_0043_ wrapper_0/_0044_ wrapper_0/_0700_ wrapper_0/_0702_ wrapper_0/_0704_
+ wrapper_0/_0410_ wrapper_0/_0412_ wrapper_0/_0738_ wrapper_0/_0739_ wrapper_0/_0143_
+ wrapper_0/_0267_ wrapper_0/_0269_ wrapper_0/_0271_ wrapper_0/_0273_ wrapper_0/clknet_4_12_0_clk_in
+ wrapper_0/clknet_4_13_0_clk_in wrapper_0/_0144_ wrapper_0/d2.r_reg\[12\] wrapper_0/d2.r_reg\[13\]
+ wrapper_0/d2.r_reg\[14\] wrapper_0/d2.r_reg\[16\] wrapper_0/d2.r_reg\[18\] wrapper_0/_0034_
+ wrapper_0/_0773_ wrapper_0/_0175_ wrapper_0/_0176_ wrapper_0/_0617_ wrapper_0/_0177_
+ wrapper_0/_0853_ wrapper_0/d2.r_reg\[50\] wrapper_0/d2.t_load\[10\] wrapper_0/d2.t_load\[11\]
+ wrapper_0/_0304_ wrapper_0/d2.t_load\[15\] wrapper_0/d2.t_load\[16\] wrapper_0/d2.t_load\[17\]
+ wrapper_0/_0372_ wrapper_0/_0373_ wrapper_0/_0374_ wrapper_0/_0375_ wrapper_0/_0376_
+ wrapper_0/_0377_ wrapper_0/_0378_ wrapper_0/_0379_ wrapper_0/_0178_ wrapper_0/_0889_
+ wrapper_0/d2.t_load\[50\] wrapper_0/d2.t_load\[51\] wrapper_0/_0890_ wrapper_0/_0891_
+ wrapper_0/_0894_ wrapper_0/_0897_ wrapper_0/_0040_ wrapper_0/_0138_ wrapper_0/_0139_
+ wrapper_0/_0140_ wrapper_0/_0690_ wrapper_0/_0692_ wrapper_0/_0694_ wrapper_0/_0695_
+ wrapper_0/_0696_ wrapper_0/_0697_ wrapper_0/_0698_ wrapper_0/_0950_ wrapper_0/_0952_
+ wrapper_0/_0953_ wrapper_0/_0956_ wrapper_0/_0957_ wrapper_0/_0958_ wrapper_0/_0959_
+ wrapper_0/_0960_ wrapper_0/_0962_ wrapper_0/_0965_ wrapper_0/_0968_ wrapper_0/clknet_0_ref_in
+ wrapper_0/clknet_1_1__leaf_ref_in wrapper_0/_0509_ wrapper_0/_0510_ wrapper_0/_0513_
+ wrapper_0/_0797_ wrapper_0/_0514_ wrapper_0/_0799_ wrapper_0/_0515_ wrapper_0/_0516_
+ wrapper_0/_0518_ wrapper_0/_0118_ wrapper_0/_0120_ wrapper_0/_0141_ wrapper_0/_0457_
+ wrapper_0/_0459_ wrapper_0/_0462_ wrapper_0/_0121_ wrapper_0/_0124_ wrapper_0/_0223_
+ wrapper_0/_0000_ wrapper_0/_0354_ wrapper_0/_0355_ wrapper_0/_0356_ wrapper_0/d2.t_load\[18\]
+ wrapper_0/_0472_ wrapper_0/_0358_ wrapper_0/_0474_ wrapper_0/_0475_ wrapper_0/_0476_
+ wrapper_0/_0477_ wrapper_0/_0478_ wrapper_0/_0359_ wrapper_0/_0482_ wrapper_0/_0485_
+ wrapper_0/_0486_ wrapper_0/_0487_ wrapper_0/d5.fll_core.corner_tmp\[0\] wrapper_0/d5.fll_core.corner_tmp\[2\]
+ wrapper_0/_0488_ wrapper_0/_0489_ wrapper_0/_0490_ wrapper_0/_0491_ wrapper_0/_0492_
+ wrapper_0/_0495_ wrapper_0/_0496_ wrapper_0/_0498_ wrapper_0/_0502_ wrapper_0/d5.fll_core.tmp\[0\]
+ wrapper_0/d5.fll_core.tmp\[1\] wrapper_0/d5.fll_core.tmp\[3\] wrapper_0/d5.fll_core.tmp\[6\]
+ wrapper_0/_0504_ wrapper_0/net43 wrapper_0/_0506_ wrapper_0/_0508_ wrapper_0/_0945_
+ wrapper_0/_0947_ wrapper_0/_0948_ wrapper_0/_0748_ wrapper_0/_0749_ wrapper_0/_0750_
+ wrapper_0/_0777_ wrapper_0/_0789_ wrapper_0/_0859_ wrapper_0/_0865_ wrapper_0/_0866_
+ wrapper_0/_0871_ wrapper_0/_0872_ wrapper_0/_0873_ wrapper_0/_0874_ wrapper_0/_0876_
+ wrapper_0/_0877_ wrapper_0/_0156_ wrapper_0/_0880_ wrapper_0/_0159_ wrapper_0/_0286_
+ wrapper_0/_0287_ wrapper_0/_0288_ wrapper_0/_0289_ wrapper_0/_0290_ wrapper_0/_0291_
+ wrapper_0/_0640_ wrapper_0/_0642_ wrapper_0/clknet_4_11_0_clk_in wrapper_0/_0644_
+ wrapper_0/_0650_ wrapper_0/_0651_ wrapper_0/_0653_ wrapper_0/_0654_ wrapper_0/_0655_
+ wrapper_0/_0657_ wrapper_0/_0658_ wrapper_0/_0661_ wrapper_0/d2.r_reg\[29\] wrapper_0/d2.r_reg\[30\]
+ wrapper_0/_0662_ wrapper_0/d2.r_reg\[32\] wrapper_0/d2.r_reg\[33\] wrapper_0/d2.r_reg\[34\]
+ wrapper_0/d2.r_reg\[36\] wrapper_0/d2.r_reg\[37\] wrapper_0/d2.r_reg\[41\] wrapper_0/_0663_
+ wrapper_0/_0664_ wrapper_0/_0665_ wrapper_0/_0666_ wrapper_0/_0669_ wrapper_0/_0670_
+ vdd wrapper_0/_0049_ wrapper_0/_0050_ wrapper_0/_0051_ wrapper_0/d2.t_load\[29\]
+ wrapper_0/_0052_ wrapper_0/d2.t_load\[33\] wrapper_0/d2.t_load\[34\] wrapper_0/d2.t_load\[39\]
+ wrapper_0/d2.t_load\[44\] wrapper_0/_0390_ wrapper_0/_0391_ wrapper_0/_0393_ wrapper_0/_0394_
+ wrapper_0/_0396_ wrapper_0/_0400_ wrapper_0/_0401_ wrapper_0/_0402_ wrapper_0/_0060_
+ wrapper_0/net12 wrapper_0/_0743_ wrapper_0/_0164_ wrapper_0/_0168_ wrapper_0/_0630_
+ wrapper_0/_0637_ wrapper_0/_0864_ wrapper_0/_0059_ wrapper_0/_0641_ wrapper_0/_0862_
+ wrapper_0/d2.t_load\[36\] wrapper_0/d2.t_load\[37\] wrapper_0/_0643_ wrapper_0/d2.t_load\[41\]
+ wrapper_0/_0863_ wrapper_0/_0868_ wrapper_0/_0645_ wrapper_0/d2.r_reg\[38\] wrapper_0/_0646_
+ wrapper_0/d2.r_reg\[42\] wrapper_0/_0647_ wrapper_0/_0649_ wrapper_0/_0292_ wrapper_0/_0403_
+ wrapper_0/_0293_ wrapper_0/_0295_ wrapper_0/_0297_ wrapper_0/net17 wrapper_0/net19
+ wrapper_0/_0061_ wrapper_0/_0163_ wrapper_0/_0744_ wrapper_0/net8 wrapper_0/net9
+ wrapper_0/_0745_ wrapper_0/_0066_ wrapper_0/_0593_ wrapper_0/d2.t_load\[43\] wrapper_0/d2.r_reg\[44\]
+ wrapper_0/_0595_ wrapper_0/d2.r_reg\[61\] wrapper_0/d2.t_load\[62\] wrapper_0/d2.r_reg\[62\]
+ wrapper_0/_0598_ wrapper_0/_0629_ wrapper_0/_0840_ wrapper_0/_0635_ wrapper_0/_0636_
+ wrapper_0/_0083_ wrapper_0/_0404_ wrapper_0/_0405_ wrapper_0/_0841_ wrapper_0/_0296_
+ wrapper_0/_0065_ wrapper_0/_0187_ wrapper_0/_0189_ wrapper_0/_0424_ wrapper_0/net26
+ wrapper_0/net27 wrapper_0/clknet_4_10_0_clk_in wrapper_0/_0315_ wrapper_0/_0316_
+ wrapper_0/_0317_ wrapper_0/_0062_ wrapper_0/clknet_4_8_0_clk_in wrapper_0/_0302_
+ wrapper_0/_0303_ wrapper_0/_0071_ wrapper_0/_0312_ wrapper_0/_0313_ wrapper_0/_0183_
+ wrapper_0/_0184_ wrapper_0/_0186_ wrapper_0/_0855_ wrapper_0/_0420_ wrapper_0/_0190_
+ wrapper_0/_0248_ wrapper_0/_0249_ wrapper_0/_0418_ wrapper_0/_0171_ wrapper_0/_0174_
+ wrapper_0/_0172_ wrapper_0/_0586_ wrapper_0/_0790_ wrapper_0/_0791_ wrapper_0/_0250_
+ wrapper_0/_0602_ wrapper_0/d2.t_load\[45\] wrapper_0/d2.t_load\[46\] wrapper_0/_0604_
+ wrapper_0/_0605_ wrapper_0/d2.t_load\[57\] wrapper_0/d2.t_load\[58\] wrapper_0/d2.t_load\[60\]
+ wrapper_0/_0173_ wrapper_0/_0618_ wrapper_0/_0620_ wrapper_0/_0622_ wrapper_0/_0624_
+ wrapper_0/_0626_ wrapper_0/_0628_ wrapper_0/_0079_ wrapper_0/_0245_ wrapper_0/_0631_
+ wrapper_0/_0406_ wrapper_0/_0409_ wrapper_0/d5.fll_core.strobe wrapper_0/d2.r_reg\[45\]
+ wrapper_0/_0733_ wrapper_0/_0734_ wrapper_0/_0735_ wrapper_0/d5.mux01.out\[3\] wrapper_0/d5.mux01.out\[5\]
+ wrapper_0/d5.mux01.out\[6\] wrapper_0/d5.mux01.out\[7\] wrapper_0/d2.r_reg\[46\]
+ wrapper_0/d2.r_reg\[47\] wrapper_0/_0736_ wrapper_0/d2.r_reg\[48\] wrapper_0/d2.r_reg\[49\]
+ wrapper_0/_0633_ wrapper_0/d2.r_reg\[51\] wrapper_0/d2.r_reg\[58\] wrapper_0/_0737_
+ wrapper_0/_0069_ wrapper_0/_0417_ wrapper_0/_0740_ wrapper_0/_0070_ wrapper_0/_0246_
+ wrapper_0/_0247_ wrapper_0/_0843_ wrapper_0/_0300_ wrapper_0/_0201_ wrapper_0/_0202_
+ wrapper_0/_0741_ wrapper_0/_0742_ wrapper_0/_0077_ wrapper_0/_0588_ wrapper_0/_0589_
+ wrapper_0/_0308_ wrapper_0/d2.r_reg\[54\] wrapper_0/d2.r_reg\[55\] wrapper_0/d2.r_reg\[56\]
+ wrapper_0/_0310_ wrapper_0/_0075_ wrapper_0/d2.r_reg\[66\] wrapper_0/d2.r_reg\[75\]
+ wrapper_0/_0836_ wrapper_0/_0838_ wrapper_0/_0414_ wrapper_0/_0415_ wrapper_0/_0076_
+ wrapper_0/_0847_ wrapper_0/_0849_ wrapper_0/_0850_ wrapper_0/_0851_ wrapper_0/_0606_
+ wrapper_0/_0607_ wrapper_0/_0608_ wrapper_0/_0609_ wrapper_0/_0611_ wrapper_0/_0086_
+ wrapper_0/_0425_ wrapper_0/d2.t_load\[54\] wrapper_0/d2.t_load\[55\] wrapper_0/d2.t_load\[65\]
+ wrapper_0/_0435_ wrapper_0/_0436_ wrapper_0/_0320_ wrapper_0/d5.fll_core.tmp\[9\]
+ wrapper_0/_0892_ wrapper_0/d5.mux01.out\[9\] wrapper_0/_0253_ wrapper_0/_0181_ wrapper_0/_0182_
+ wrapper_0/_0095_ wrapper_0/_0096_ wrapper_0/_0192_ wrapper_0/_0584_ wrapper_0/_0585_
+ wrapper_0/_0781_ wrapper_0/_0782_ wrapper_0/clknet_4_2_0_clk_in wrapper_0/clknet_4_3_0_clk_in
+ wrapper_0/_0195_ wrapper_0/_0590_ wrapper_0/_0592_ wrapper_0/_0792_ wrapper_0/_0200_
+ wrapper_0/_0594_ wrapper_0/_0084_ wrapper_0/_0085_ wrapper_0/_0568_ wrapper_0/_0569_
+ wrapper_0/_0570_ wrapper_0/_0571_ wrapper_0/_0427_ wrapper_0/_0429_ wrapper_0/_0572_
+ wrapper_0/_0434_ wrapper_0/d2.r_reg\[63\] wrapper_0/_0579_ wrapper_0/_0318_ wrapper_0/_0319_
+ wrapper_0/d2.r_reg\[68\] wrapper_0/_0321_ wrapper_0/_0323_ wrapper_0/_0324_ wrapper_0/d2.r_reg\[72\]
+ wrapper_0/_0581_ wrapper_0/_0087_ wrapper_0/_0825_ wrapper_0/_0088_ wrapper_0/_0089_
+ wrapper_0/_0828_ wrapper_0/_0094_ wrapper_0/net23 wrapper_0/net24 wrapper_0/net25
+ wrapper_0/_0833_ wrapper_0/_0834_ wrapper_0/_0582_ wrapper_0/_0583_ wrapper_0/_0839_
+ wrapper_0/_0193_ wrapper_0/_0194_ wrapper_0/_0196_ wrapper_0/_0433_ wrapper_0/_0564_
+ wrapper_0/_0091_ wrapper_0/_0092_ wrapper_0/_0197_ wrapper_0/_0576_ wrapper_0/net20
+ wrapper_0/net21 wrapper_0/net22 wrapper_0/_0829_ wrapper_0/_0830_ wrapper_0/_0831_
+ wrapper_0/_0832_ wrapper_0/_0577_ wrapper_0/_0578_ wrapper_0/_0330_ wrapper_0/d2.r_reg\[70\]
+ wrapper_0/_0431_ wrapper_0/_0432_ wrapper_0/_0559_ wrapper_0/_0560_ wrapper_0/_0561_
+ wrapper_0/_0441_ wrapper_0/_0442_ wrapper_0/_0562_ wrapper_0/clknet_4_1_0_clk_in
+ wrapper_0/_0203_ wrapper_0/_0204_ wrapper_0/_0563_ wrapper_0/_0205_ wrapper_0/_0566_
+ wrapper_0/_0331_ wrapper_0/_0332_ wrapper_0/_0333_ wrapper_0/_0793_ wrapper_0/_0207_
+ wrapper_0/_0334_ wrapper_0/_0337_ wrapper_0/_0104_ wrapper_0/_0547_ wrapper_0/_0548_
+ wrapper_0/_0549_ wrapper_0/_0550_ wrapper_0/_0551_ wrapper_0/_0817_ wrapper_0/_0575_
+ wrapper_0/_0552_ wrapper_0/_0553_ wrapper_0/_0554_ wrapper_0/_0555_ wrapper_0/_0556_
+ wrapper_0/d2.r_reg\[77\] wrapper_0/d2.r_reg\[79\] wrapper_0/d2.r_reg\[81\] wrapper_0/net30
+ wrapper_0/net31 wrapper_0/net32 wrapper_0/net33 wrapper_0/_0819_ wrapper_0/_0821_
+ wrapper_0/_0098_ wrapper_0/_0100_ wrapper_0/_0101_ wrapper_0/_0102_ wrapper_0/_0824_
+ wrapper_0/clknet_4_0_0_clk_in wrapper_0/_0557_ wrapper_0/_0453_ wrapper_0/_0460_
+ wrapper_0/_0973_ wrapper_0/_0974_ wrapper_0/_0976_ wrapper_0/_0977_ wrapper_0/_0980_
+ wrapper_0/_0981_ wrapper_0/_0984_ wrapper_0/_0985_ wrapper_0/_0986_ wrapper_0/_0990_
+ wrapper_0/_0991_ wrapper_0/_0461_ wrapper_0/_0761_ wrapper_0/_0762_ wrapper_0/_0763_
+ wrapper_0/_0764_ wrapper_0/_0765_ wrapper_0/_0766_ wrapper_0/_0768_ wrapper_0/_0769_
+ wrapper_0/_0785_ wrapper_0/_0016_ wrapper_0/_0011_ wrapper_0/_0500_ wrapper_0/_0501_
+ wrapper_0/_0112_ wrapper_0/_0528_ wrapper_0/_0529_ wrapper_0/_0532_ wrapper_0/_0012_
+ wrapper_0/_0013_ wrapper_0/_0123_ wrapper_0/_0015_ wrapper_0/_0128_ wrapper_0/_0236_
+ wrapper_0/_0237_ wrapper_0/_0240_ wrapper_0/d5.fll_core.counter2.count\[1\] wrapper_0/d5.fll_core.counter2.count\[2\]
+ wrapper_0/d5.fll_core.counter2.count\[5\] wrapper_0/d5.fll_core.counter2.count\[6\]
+ wrapper_0/d5.fll_core.counter2.count\[7\] wrapper_0/d5.fll_core.counter2.count\[8\]
+ wrapper_0/_0243_ wrapper_0/_0244_ wrapper_0/_0908_ wrapper_0/net42 wrapper_0/_0136_
+ wrapper_0/_0137_ wrapper_0/_0848_ wrapper_0/_0264_ wrapper_0/_0365_ wrapper_0/d2.t_load\[3\]
+ wrapper_0/clknet_4_6_0_clk_in wrapper_0/d2.t_load\[4\] wrapper_0/d2.t_load\[7\]
+ wrapper_0/d2.t_load\[8\] wrapper_0/d2.t_load\[9\] wrapper_0/_0306_ wrapper_0/_0786_
+ wrapper_0/_0366_ wrapper_0/_0367_ wrapper_0/_0368_ wrapper_0/clknet_4_7_0_clk_in
+ wrapper_0/_0616_ wrapper_0/_0025_ wrapper_0/_0026_ wrapper_0/_0030_ wrapper_0/_0260_
+ wrapper_0/_0073_ wrapper_0/d2.r_reg\[4\] wrapper_0/d2.r_reg\[5\] wrapper_0/d2.r_reg\[6\]
+ wrapper_0/d2.r_reg\[7\] wrapper_0/d2.r_reg\[10\] wrapper_0/_0129_ wrapper_0/_0899_
+ wrapper_0/_0901_ wrapper_0/_0904_ wrapper_0/d5.fll_core.tmp\[8\] wrapper_0/_0905_
+ wrapper_0/_0259_ wrapper_0/_0130_ wrapper_0/d5.mux01.out\[8\] wrapper_0/_0131_ wrapper_0/_0179_
+ wrapper_0/_0706_ wrapper_0/_0708_ wrapper_0/_0709_ wrapper_0/_0710_ wrapper_0/_0711_
+ wrapper_0/_0712_ wrapper_0/_0713_ wrapper_0/_0714_ wrapper_0/_0715_ wrapper_0/_0716_
+ wrapper_0/_0717_ wrapper_0/_0718_ wrapper_0/_0719_ wrapper_0/_0720_ wrapper_0/_0721_
+ wrapper_0/_0722_ wrapper_0/_0263_ wrapper_0/_0134_ wrapper_0/_0074_ wrapper_0/d2.t_load\[1\]
+ wrapper_0/_0814_ wrapper_0/_0530_ wrapper_0/_0815_ wrapper_0/_0774_ wrapper_0/_0541_
+ wrapper_0/_0542_ wrapper_0/_0543_ wrapper_0/_0544_ wrapper_0/_0545_ wrapper_0/_0546_
+ wrapper_0/_0221_ wrapper_0/_0816_ wrapper_0/_0105_ wrapper_0/net1 wrapper_0/_0106_
+ wrapper_0/_0349_ wrapper_0/d2.r_reg\[84\] wrapper_0/net2 wrapper_0/d2.r_reg\[85\]
+ wrapper_0/_0256_ wrapper_0/_0023_ wrapper_0/_0802_ wrapper_0/_0115_ wrapper_0/_0783_
+ wrapper_0/_0803_ wrapper_0/_0211_ wrapper_0/net28 wrapper_0/_0212_ wrapper_0/_0220_
+ wrapper_0/_0519_ wrapper_0/_0723_ wrapper_0/net36 wrapper_0/_0805_ wrapper_0/_0725_
+ wrapper_0/_0524_ wrapper_0/_0806_ wrapper_0/_0794_ wrapper_0/_0255_ wrapper_0/_0340_
+ wrapper_0/_0116_ wrapper_0/_0809_ wrapper_0/_0810_ wrapper_0/_0450_ wrapper_0/_0811_
+ wrapper_0/_0214_ wrapper_0/_0216_ wrapper_0/_0812_ wrapper_0/_0813_ wrapper_0/_0344_
+ wrapper_0/_0521_ wrapper_0/_0522_ wrapper_0/_0362_ wrapper_0/_0525_ wrapper_0/_0526_
+ wrapper_0/_0527_ wrapper_0/_0909_ wrapper_0/_0910_ wrapper_0/_0795_ wrapper_0/_0345_
+ wrapper_0/_0347_ wrapper_0/_0348_ wrapper_0/_0108_ wrapper_0/_0533_ wrapper_0/_0534_
+ wrapper_0/_0536_ wrapper_0/net16 wrapper_0/_0109_ wrapper_0/_0537_ wrapper_0/_0540_
+ wrapper_0/_0451_ wrapper_0/_0111_ wrapper_0/_0350_ wrapper_0/_0449_ wrapper_0/d2.r_reg\[86\]
+ wrapper_0/d2.r_reg\[87\] wrapper_0/d2.r_reg\[88\] wrapper_0/d2.r_reg\[89\] wrapper_0/d2.r_reg\[90\]
+ wrapper_0/d2.t_load\[93\] wrapper_0/d2.t_load\[94\] wrapper_0/d2.r_reg\[93\] wrapper_0/d2.r_reg\[95\]
+ wrapper_0/d2.t_load\[0\] wrapper_0/net39 wrapper_0/net4 wrapper_0/net40 wrapper_0/_0456_
+ wrapper_0/_0804_ wrapper_0/_0728_ wrapper_0/_0342_ wrapper_0/_0127_ wrapper_0/_0113_
+ wrapper_0/_0114_ wrapper_0/_0343_ wrapper_0/_0447_ wrapper_0/_0448_ full_vco_1_0/b0
+ full_vco_1_0/b1 full_vco_1_0/b2 slopebuf_0/bit0 slopebuf_0/bit1 slopebuf_0/bit2
+ r2r_8_1/b0 r2r_8_1/b1 r2r_8_1/b2 r2r_8_1/b3 r2r_8_1/b4 r2r_8_1/b5 r2r_8_1/b6 r2r_8_1/b7
+ r2r_8_0/b0 r2r_8_0/b1 r2r_8_0/b2 r2r_8_0/b3 r2r_8_0/b4 r2r_8_0/b5 r2r_8_0/b6 r2r_8_0/b7
+ wrapper_0/_0003_ wrapper_0/_0004_ wrapper_0/_0005_ wrapper_0/_0007_ wrapper_0/_0008_
+ wrapper_0/_0009_ wrapper_0/_0228_ wrapper_0/_0231_ wrapper_0/_0232_ wrapper_0/_0233_
+ wrapper_0/_0234_ wrapper_0/_0458_ wrapper_0/_0731_ wrapper_0/_0756_ wrapper_0/_0758_
+ wrapper_0/_0759_ wrapper_0/_0911_ wrapper_0/_0916_ wrapper_0/_0917_ wrapper_0/_0935_
+ wrapper_0/clknet_0_vco_in wrapper_0/clknet_1_0__leaf_vco_in wrapper_0/clknet_1_1__leaf_vco_in
+ wrapper_0/d5.fll_core.corner_tmp\[1\] wrapper_0/d5.fll_core.counter1.count\[9\]
+ wrapper_0/net5 wrapper_0/_0682_ wrapper_0/_0687_ wrapper_0/_0688_ wrapper_0/_0157_
+ wrapper_0/_0041_ wrapper_0/_0046_ wrapper_0/_0047_ wrapper_0/_0776_ wrapper_0/_0879_
+ wrapper_0/_0887_ wrapper_0/_0152_ wrapper_0/_0153_ wrapper_0/_0279_ wrapper_0/_0922_
+ wrapper_0/_0924_ wrapper_0/_0926_ wrapper_0/_0928_ wrapper_0/_0929_ wrapper_0/_0933_
+ wrapper_0/_0280_ wrapper_0/clknet_0_clk_in wrapper_0/_0281_ wrapper_0/_0380_ wrapper_0/_0382_
+ wrapper_0/_0385_ wrapper_0/_0386_ wrapper_0/_0392_ wrapper_0/d2.r_reg\[19\] wrapper_0/d2.r_reg\[20\]
+ wrapper_0/d2.r_reg\[23\] wrapper_0/d2.r_reg\[26\] wrapper_0/d2.t_load\[12\] wrapper_0/d2.t_load\[22\]
+ wrapper_0/d2.t_load\[26\] wrapper_0/_0155_ wrapper_0/d5.fll_core.counter1.count\[3\]
+ wrapper_0/_0466_ wrapper_0/_0676_ wrapper_0/_0680_ wrapper_0/_0033_ wrapper_0/_0142_
+ wrapper_0/_0625_ wrapper_0/_0268_ wrapper_0/_0270_ wrapper_0/_0272_ wrapper_0/_0274_
+ wrapper_0/_0145_ wrapper_0/_0691_ wrapper_0/_0693_ wrapper_0/_0699_ wrapper_0/_0701_
+ wrapper_0/_0703_ wrapper_0/_0705_ wrapper_0/_0707_ wrapper_0/_0035_ wrapper_0/d2.r_reg\[11\]
+ wrapper_0/d2.r_reg\[15\] wrapper_0/d2.r_reg\[17\] wrapper_0/_0036_ wrapper_0/_0037_
+ wrapper_0/_0038_ wrapper_0/_0775_ wrapper_0/d2.r_reg\[52\] wrapper_0/_0039_ wrapper_0/_0854_
+ wrapper_0/_0031_ wrapper_0/d2.t_load\[49\] wrapper_0/_0032_ wrapper_0/_0895_ wrapper_0/_0896_
+ wrapper_0/_0898_ wrapper_0/_0411_ wrapper_0/_0483_ wrapper_0/_0944_ wrapper_0/_0946_
+ wrapper_0/_0949_ wrapper_0/_0951_ wrapper_0/_0954_ wrapper_0/_0955_ wrapper_0/_0961_
+ wrapper_0/_0963_ wrapper_0/_0964_ wrapper_0/_0966_ wrapper_0/_0967_ wrapper_0/_0969_
+ wrapper_0/_0970_ wrapper_0/_0971_ wrapper_0/_0484_ wrapper_0/_0493_ wrapper_0/clknet_1_0__leaf_ref_in
+ wrapper_0/_0494_ wrapper_0/_0497_ wrapper_0/_0499_ wrapper_0/_0503_ wrapper_0/_0505_
+ wrapper_0/_0784_ wrapper_0/_0796_ wrapper_0/_0507_ wrapper_0/_0511_ wrapper_0/_0512_
+ wrapper_0/_0517_ wrapper_0/_0117_ wrapper_0/_0119_ wrapper_0/_0224_ wrapper_0/d2.t_load\[14\]
+ wrapper_0/_0122_ wrapper_0/_0125_ wrapper_0/_0351_ wrapper_0/_0352_ wrapper_0/_0353_
+ wrapper_0/_0471_ wrapper_0/d5.fll_core.tmp\[2\] wrapper_0/d5.fll_core.tmp\[4\] wrapper_0/d5.fll_core.tmp\[5\]
+ wrapper_0/d5.fll_core.tmp\[7\] wrapper_0/_0479_ wrapper_0/_0481_ wrapper_0/_0747_
+ wrapper_0/_0160_ wrapper_0/_0161_ wrapper_0/_0162_ wrapper_0/_0387_ wrapper_0/_0166_
+ wrapper_0/_0395_ wrapper_0/_0167_ wrapper_0/_0048_ wrapper_0/_0053_ wrapper_0/_0054_
+ wrapper_0/_0055_ wrapper_0/_0056_ wrapper_0/clknet_4_14_0_clk_in wrapper_0/_0057_
+ wrapper_0/_0627_ wrapper_0/_0656_ wrapper_0/_0659_ wrapper_0/d2.r_reg\[35\] wrapper_0/d2.r_reg\[39\]
+ wrapper_0/d2.r_reg\[40\] wrapper_0/_0660_ wrapper_0/_0667_ wrapper_0/_0668_ wrapper_0/_0283_
+ wrapper_0/d2.t_load\[32\] wrapper_0/d2.t_load\[35\] wrapper_0/d2.t_load\[40\] wrapper_0/_0284_
+ wrapper_0/d2.t_load\[56\] wrapper_0/_0285_ wrapper_0/_0294_ wrapper_0/net13 wrapper_0/net14
+ wrapper_0/net15 wrapper_0/_0638_ wrapper_0/_0639_ wrapper_0/_0648_ wrapper_0/d2.t_load\[38\]
+ wrapper_0/_0746_ wrapper_0/d2.t_load\[42\] wrapper_0/_0397_ wrapper_0/_0867_ wrapper_0/_0869_
+ wrapper_0/_0398_ wrapper_0/d2.r_reg\[43\] wrapper_0/_0399_ wrapper_0/net10 wrapper_0/net11
+ wrapper_0/_0165_ wrapper_0/_0169_ wrapper_0/_0058_ wrapper_0/_0063_ wrapper_0/_0423_
+ wrapper_0/d2.t_load\[61\] wrapper_0/_0596_ wrapper_0/_0597_ wrapper_0/_0298_ wrapper_0/_0299_
+ wrapper_0/_0599_ wrapper_0/d2.r_reg\[60\] wrapper_0/_0861_ wrapper_0/_0170_ wrapper_0/_0188_
+ wrapper_0/_0634_ wrapper_0/_0081_ wrapper_0/_0082_ wrapper_0/_0842_ wrapper_0/_0778_
+ wrapper_0/net18 wrapper_0/_0421_ wrapper_0/_0422_ wrapper_0/_0064_ wrapper_0/_0846_
+ wrapper_0/_0600_ wrapper_0/_0601_ wrapper_0/_0603_ wrapper_0/_0619_ wrapper_0/_0621_
+ wrapper_0/_0185_ wrapper_0/d2.t_load\[47\] wrapper_0/d2.t_load\[48\] wrapper_0/clknet_4_9_0_clk_in
+ wrapper_0/_0623_ wrapper_0/d2.t_load\[59\] wrapper_0/_0779_ wrapper_0/d2.t_load\[63\]
+ wrapper_0/_0068_ wrapper_0/_0632_ wrapper_0/_0072_ wrapper_0/_0078_ wrapper_0/_0301_
+ wrapper_0/_0305_ wrapper_0/_0314_ wrapper_0/d5.mux01.out\[0\] wrapper_0/d5.mux01.out\[1\]
+ wrapper_0/d5.mux01.out\[2\] wrapper_0/d5.mux01.out\[4\] wrapper_0/_0080_ wrapper_0/_0856_
+ wrapper_0/_0407_ wrapper_0/_0251_ wrapper_0/_0252_ wrapper_0/_0408_ wrapper_0/_0857_
+ wrapper_0/_0419_ wrapper_0/_0858_ wrapper_0/d2.r_reg\[57\] wrapper_0/d2.r_reg\[59\]
+ wrapper_0/_0860_ wrapper_0/_0844_ wrapper_0/_0845_ wrapper_0/_0067_ wrapper_0/_0826_
+ wrapper_0/_0827_ wrapper_0/_0835_ wrapper_0/_0837_ wrapper_0/_0311_ wrapper_0/_0206_
+ wrapper_0/_0416_ wrapper_0/_0322_ wrapper_0/_0610_ wrapper_0/_0612_ wrapper_0/_0613_
+ wrapper_0/_0614_ wrapper_0/_0325_ wrapper_0/_0326_ wrapper_0/d2.r_reg\[64\] wrapper_0/d2.r_reg\[65\]
+ wrapper_0/d2.r_reg\[67\] wrapper_0/d2.r_reg\[69\] wrapper_0/d2.r_reg\[71\] wrapper_0/d2.r_reg\[73\]
+ wrapper_0/d2.r_reg\[74\] wrapper_0/d2.r_reg\[76\] wrapper_0/d2.r_reg\[78\] wrapper_0/d2.r_reg\[80\]
+ wrapper_0/d2.r_reg\[82\] wrapper_0/d2.r_reg\[83\] wrapper_0/_0327_ wrapper_0/_0426_
+ wrapper_0/_0428_ wrapper_0/_0430_ wrapper_0/_0437_ wrapper_0/_0438_ wrapper_0/_0439_
+ wrapper_0/_0440_ wrapper_0/_0443_ wrapper_0/_0444_ wrapper_0/_0328_ wrapper_0/_0329_
+ wrapper_0/_0335_ wrapper_0/_0336_ wrapper_0/_0338_ wrapper_0/_0208_ wrapper_0/d2.t_load\[64\]
+ wrapper_0/_0209_ wrapper_0/_0210_ wrapper_0/_0090_ wrapper_0/_0093_ wrapper_0/_0097_
+ wrapper_0/_0180_ wrapper_0/_0099_ wrapper_0/_0103_ wrapper_0/_0191_ wrapper_0/_0198_
+ wrapper_0/_0254_ wrapper_0/_0558_ wrapper_0/_0565_ wrapper_0/_0567_ wrapper_0/_0573_
+ wrapper_0/_0574_ wrapper_0/_0580_ wrapper_0/_0587_ wrapper_0/_0591_ wrapper_0/_0780_
+ wrapper_0/_0199_ wrapper_0/_0309_ wrapper_0/net29 wrapper_0/net34 wrapper_0/net35
+ wrapper_0/_0818_ wrapper_0/_0820_ wrapper_0/_0822_ wrapper_0/_0823_ wrapper_0/_0360_
+ wrapper_0/_0361_ wrapper_0/_0363_ wrapper_0/_0767_ wrapper_0/_0770_ wrapper_0/_0771_
+ wrapper_0/_0531_ wrapper_0/_0801_ wrapper_0/_0807_ wrapper_0/_0808_ wrapper_0/_0019_
+ wrapper_0/_0020_ wrapper_0/d2.r_reg\[91\] wrapper_0/d2.r_reg\[92\] wrapper_0/_0217_
+ wrapper_0/_0218_ wrapper_0/_0219_ wrapper_0/_0903_ wrapper_0/_0014_ wrapper_0/_0017_
+ wrapper_0/_0018_ wrapper_0/d5.fll_core.counter2.count\[0\] wrapper_0/d5.fll_core.counter2.count\[3\]
+ wrapper_0/d5.fll_core.counter2.count\[4\] wrapper_0/d5.fll_core.counter2.count\[9\]
+ wrapper_0/_0235_ wrapper_0/_0238_ wrapper_0/_0452_ wrapper_0/_0239_ wrapper_0/_0241_
+ wrapper_0/_0242_ wrapper_0/_0126_ wrapper_0/_0346_ wrapper_0/_0972_ wrapper_0/_0975_
+ wrapper_0/net41 wrapper_0/_0978_ wrapper_0/_0979_ wrapper_0/_0982_ wrapper_0/_0983_
+ wrapper_0/_0988_ wrapper_0/_0989_ wrapper_0/_0357_ wrapper_0/_0906_ wrapper_0/_0907_
+ wrapper_0/_0029_ wrapper_0/d2.t_load\[6\] wrapper_0/_0265_ wrapper_0/_0266_ wrapper_0/_0135_
+ wrapper_0/d2.r_reg\[3\] wrapper_0/_0364_ wrapper_0/_0024_ wrapper_0/_0852_ wrapper_0/_0027_
+ wrapper_0/_0028_ wrapper_0/d2.r_reg\[8\] wrapper_0/_0369_ wrapper_0/_0370_ wrapper_0/d2.r_reg\[9\]
+ wrapper_0/_0413_ wrapper_0/_0132_ wrapper_0/d2.r_reg\[53\] wrapper_0/_0133_ wrapper_0/_0724_
+ wrapper_0/_0726_ wrapper_0/_0615_ wrapper_0/d2.t_load\[2\] wrapper_0/_0371_ wrapper_0/_0261_
+ wrapper_0/_0893_ wrapper_0/_0307_ wrapper_0/_0900_ wrapper_0/_0987_ wrapper_0/d2.t_load\[52\]
+ wrapper_0/d2.t_load\[53\] wrapper_0/_0902_ wrapper_0/_0262_ wrapper_0/_0258_ wrapper_0/d2.t_load\[5\]
+ wrapper_0/_0446_ wrapper_0/_0727_ wrapper_0/net3 wrapper_0/_0772_ wrapper_0/_0454_
+ wrapper_0/_0455_ wrapper_0/d2.r_reg\[94\] wrapper_0/d2.r_reg\[2\] wrapper_0/_0107_
+ wrapper_0/clknet_4_4_0_clk_in wrapper_0/d2.r_reg\[1\] wrapper_0/_0339_ wrapper_0/_0341_
+ wrapper_0/_0729_ wrapper_0/_0021_ wrapper_0/_0022_ wrapper_0/_0257_ wrapper_0/_0445_
+ wrapper_0/_0110_ wrapper_0/d2.t_load\[95\] wrapper_0/_0213_ wrapper_0/_0535_ wrapper_0/_0538_
+ wrapper_0/_0523_ wrapper_0/_0539_ wrapper_0/_0222_ wrapper_0/clknet_4_5_0_clk_in
+ wrapper_0/_0520_ wrapper_0/net37 wrapper_0/net38 wrapper_0/_0215_ vss wrapper
Xinv_buffer2_1 ref_in wrapper_0/ref_in vdd vss inv_buffer2
Xinv_buffer2_3 inv_buffer2_3/in1 slopebuf_0/clk_in vdd vss inv_buffer2
Xinv_buffer2_2 ref_in inv_buffer2_0/in1 vdd vss inv_buffer2
Xsspd_0 sspd_0/ref_in sspd_0/vco_in sspd_0/vbias sspd_0/v_out vdd vss sspd
Xvoltage_control_0 r2r_10_0/vout sspd_0/v_out vdd full_vco_1_0/vdelay wrapper_0/lock
+ vss voltage_control
Xfull_vco_1_0 full_vco_1_0/out3 wrapper_0/vco_in r2r_8_0/vout inv_buffer2_3/in1 out
+ full_vco_1_0/b0 full_vco_1_0/b1 full_vco_1_0/b2 full_vco_1_0/vdelay vdd vss full_vco_1
.ends

.subckt Standalone_mosfet_32f signal_out signal_in gnd
X0 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
D0 gnd signal_in sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X11 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X27 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X29 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X30 signal_out signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 gnd signal_in signal_out gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt RF_switch Toggle Port3 Port1 Port2 Vdd Gnd
D0 Gnd a_n50301_32455# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X0 Vdd Toggle a_n50301_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X1 Gnd a_n50301_32455# a_3046_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X2 a_4630_15090# a_4948_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X3 a_3994_15090# a_3676_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X4 Gnd a_n50301_32455# a_3046_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X5 a_n50301_32455# Toggle Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
R0 Port3 Port2 sky130_fd_pr__res_generic_m5 w=3.47e+06u l=1.1155e+07u
X6 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X7 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X8 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X9 a_3046_32455# a_n50301_32455# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X10 Gnd a_166_n5749# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X11 a_n50301_32455# Toggle Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X12 a_3994_15090# a_4312_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X13 Gnd Toggle a_n50301_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X14 a_n47356_15090# a_n50301_32455# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X15 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X16 a_n44176_15090# a_n43858_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X17 Gnd a_166_n5749# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X18 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X19 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X20 Port1 a_n42904_n5603# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X21 a_3358_15090# a_3676_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X22 Gnd a_166_n5749# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X23 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X24 Gnd a_n42904_4445# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X25 a_3046_32455# a_n50301_32455# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X26 Gnd a_166_n5749# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X27 a_3046_32455# a_n50301_32455# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X28 Gnd Toggle a_n50301_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X29 a_n43540_15090# a_n43222_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X30 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X31 Vdd Toggle a_n50301_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X32 Port1 a_n42904_n5603# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X33 Gnd a_n42904_4445# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X34 a_2722_15090# a_3040_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X35 a_n50301_32455# Toggle Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X36 a_n47356_15090# a_n47038_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X37 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X38 Port2 a_154_4444# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X39 a_n46084_15090# a_n46402_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X40 Gnd a_166_n5749# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X41 Port2 a_154_4444# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X42 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X43 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X44 a_n43540_15090# a_n43858_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X45 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X46 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X47 a_3046_32455# a_n50301_32455# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X48 Port1 a_n42904_n5603# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X49 Gnd a_n50301_32455# a_3046_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X50 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X51 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X52 Gnd a_n50301_32455# a_3046_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X53 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X54 a_3358_15090# a_3040_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X55 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X56 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X57 Gnd a_n42904_4445# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X58 Port1 a_n42904_n5603# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X59 a_n50301_32455# Toggle Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X60 a_166_n5749# a_154_4444# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.8145e+07u
X61 a_n50301_32455# Toggle Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X62 Port2 a_154_4444# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X63 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X64 a_6538_15090# a_3046_32455# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X65 Gnd Toggle a_n50301_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X66 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X67 Port1 a_n42904_n5603# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X68 a_n46720_15090# a_n46402_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X69 Vdd a_n50301_32455# a_3046_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X70 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X71 Vdd Toggle a_n50301_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X72 a_n42904_15090# a_n43222_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X73 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X74 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X75 a_5902_15090# a_6220_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X76 Gnd a_n42904_4445# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X77 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X78 a_n50301_32455# Toggle Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X79 a_3046_32455# a_n50301_32455# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X80 a_2722_15090# a_2404_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X81 a_n46720_15090# a_n47038_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X82 a_n46084_15090# a_n45766_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X83 Gnd a_n42904_4445# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X84 Port2 a_154_4444# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X85 Port2 a_154_4444# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X86 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X87 a_6538_15090# a_6220_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X88 a_5266_15090# a_5584_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X89 a_154_4444# a_2404_15090# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=5.0495e+07u
X90 Vdd a_n50301_32455# a_3046_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X91 Gnd a_166_n5749# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X92 Vdd a_n50301_32455# a_3046_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X93 a_3046_32455# a_n50301_32455# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X94 a_n50301_32455# Toggle Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X95 a_3046_32455# a_n50301_32455# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X96 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X97 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X98 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X99 a_3046_32455# a_n50301_32455# Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X100 Port1 a_n42904_n5603# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X101 Gnd Toggle a_n50301_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X102 Gnd a_166_n5749# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X103 Port2 a_154_4444# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X104 Gnd a_166_n5749# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X105 a_2404_15090# a_2404_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X106 Vdd Toggle a_n50301_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X107 a_n45448_15090# a_n45766_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X108 a_n44812_15090# a_n44494_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X109 Port2 a_154_4444# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X110 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X111 Port1 a_n42904_n5603# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X112 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X113 a_3046_32455# a_n50301_32455# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
R1 Port1 Port3 sky130_fd_pr__res_generic_m5 w=3.47e+06u l=1.1155e+07u
X114 Gnd a_166_n5749# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X115 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X116 a_5266_15090# a_4948_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X117 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X118 a_5902_15090# a_5584_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X119 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X120 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
D1 Gnd Toggle sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06u area=2.025e+11p
X121 Vdd Toggle a_n50301_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X122 Port1 a_n42904_n5603# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X123 a_n42904_n5603# a_n42904_4445# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.808e+07u
X124 Gnd a_n42904_4445# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X125 a_n42904_4445# a_n42904_15090# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=5.0435e+07u
X126 a_n50301_32455# Toggle Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X127 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X128 a_n50301_32455# Toggle Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X129 Port2 a_166_n5749# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X130 Port2 a_154_4444# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X131 Gnd a_n42904_4445# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X132 Port1 a_n42904_n5603# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X133 a_n45448_15090# a_n45130_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X134 a_n44176_15090# a_n44494_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X135 Gnd a_n50301_32455# a_3046_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X136 a_n44812_15090# a_n45130_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X137 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X138 Gnd Toggle a_n50301_32455# Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X139 Gnd a_n42904_n5603# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X140 Gnd a_n42904_4445# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X141 Vdd a_n50301_32455# a_3046_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X142 Gnd a_n42904_4445# Port1 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X143 Vdd a_n50301_32455# a_3046_32455# Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X144 Gnd a_154_4444# Port2 Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X145 a_4630_15090# a_4312_24522# Gnd sky130_fd_pr__res_xhigh_po w=350000u l=4.5e+07u
X146 a_3046_32455# a_n50301_32455# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X147 a_n50301_32455# Toggle Vdd Vdd sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X148 Port2 a_154_4444# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X149 Port1 a_n42904_4445# Gnd Gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_16 VGND VPWR Y A VNB VPB
X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X11 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X25 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X26 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X32 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X33 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X35 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X37 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_4 VPWR VGND A Y VNB VPB
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_2 VPWR VGND Y A VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_sc_hd__clkinv_8 VGND VPWR Y A VNB VPB
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
.ends

.subckt out_buf in out vdd vss
Xsky130_fd_sc_hd__clkinv_16_0 vss vdd out sky130_fd_sc_hd__clkinv_16_5/Y vss vdd sky130_fd_sc_hd__clkinv_16
Xsky130_fd_sc_hd__clkinv_16_1 vss vdd out sky130_fd_sc_hd__clkinv_16_5/Y vss vdd sky130_fd_sc_hd__clkinv_16
Xsky130_fd_sc_hd__clkinv_16_2 vss vdd out sky130_fd_sc_hd__clkinv_16_5/Y vss vdd sky130_fd_sc_hd__clkinv_16
Xsky130_fd_sc_hd__clkinv_4_0 vdd vss sky130_fd_sc_hd__clkinv_4_0/A sky130_fd_sc_hd__clkinv_8_0/A
+ vss vdd sky130_fd_sc_hd__clkinv_4
Xsky130_fd_sc_hd__clkinv_16_3 vss vdd out sky130_fd_sc_hd__clkinv_16_5/Y vss vdd sky130_fd_sc_hd__clkinv_16
Xsky130_fd_sc_hd__clkinv_16_4 vss vdd sky130_fd_sc_hd__clkinv_16_5/Y sky130_fd_sc_hd__clkinv_16_6/Y
+ vss vdd sky130_fd_sc_hd__clkinv_16
Xsky130_fd_sc_hd__clkinv_16_5 vss vdd sky130_fd_sc_hd__clkinv_16_5/Y sky130_fd_sc_hd__clkinv_16_6/Y
+ vss vdd sky130_fd_sc_hd__clkinv_16
Xsky130_fd_sc_hd__clkinv_16_6 vss vdd sky130_fd_sc_hd__clkinv_16_6/Y sky130_fd_sc_hd__clkinv_8_0/Y
+ vss vdd sky130_fd_sc_hd__clkinv_16
Xsky130_fd_sc_hd__clkinv_2_0 vdd vss sky130_fd_sc_hd__clkinv_4_0/A in vss vdd sky130_fd_sc_hd__clkinv_2
Xsky130_fd_sc_hd__clkinv_8_0 vss vdd sky130_fd_sc_hd__clkinv_8_0/Y sky130_fd_sc_hd__clkinv_8_0/A
+ vss vdd sky130_fd_sc_hd__clkinv_8
.ends

.subckt Standalone_mosfet_150f signal_in signal_out gnd
X0 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X1 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X11 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X13 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X15 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X19 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X21 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X22 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X23 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X24 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X25 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X26 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X27 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X28 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X29 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X30 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X31 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X32 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X33 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X34 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X35 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X36 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X37 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X38 a_n823_n13264# gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X39 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X40 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X41 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X42 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X43 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X44 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X45 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X46 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X47 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X48 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X49 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X50 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X51 gnd gnd a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X52 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X53 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X54 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X55 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X56 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X57 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X58 gnd gnd a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X59 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X60 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X61 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X62 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X63 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X64 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X65 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X66 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X67 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X68 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X69 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X70 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X71 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X72 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X73 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X74 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X75 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X76 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X77 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X78 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X79 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X80 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X81 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X82 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X83 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X84 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X85 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X86 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X87 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X88 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X89 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X90 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X91 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X92 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X93 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X94 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X95 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X96 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X97 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X98 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X99 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X100 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X101 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X102 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X103 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X104 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X105 a_5019_n13264# gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X106 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X107 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X108 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X109 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X110 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X111 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X112 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X113 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X114 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X115 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X116 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X117 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X118 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X119 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X120 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X121 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X122 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X123 a_n1709_n16448# gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X124 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X125 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X126 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X127 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X128 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X129 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X130 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X131 gnd gnd a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X132 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X133 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X134 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X135 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X136 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X137 a_5115_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X138 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X139 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X140 a_n727_n17334# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X141 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X142 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X143 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X144 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X145 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X146 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X147 gnd signal_in a_8203_n16352# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X148 a_5019_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X149 gnd gnd gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X150 gnd signal_in a_n823_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X151 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X152 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X153 gnd signal_in a_5115_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X154 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X155 gnd signal_in a_n727_n17334# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X156 a_n1709_n16448# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X157 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X158 gnd signal_in a_n1709_n16448# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X159 a_n823_n13264# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X160 a_8203_n16352# signal_in gnd gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X161 gnd signal_in a_5019_n13264# gnd sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
.ends

.subckt user_analog_project_wrapper wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10]
+ wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16]
+ wbs_adr_i[17] wbs_adr_i[1] wbs_adr_i[2] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[1]
+ wbs_dat_i[2] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[1] wbs_dat_o[2] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i wbs_dat_i[17] wbs_dat_i[18]
+ wbs_dat_i[19] wbs_adr_i[18] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23]
+ wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29]
+ wbs_adr_i[19] wbs_dat_i[30] wbs_dat_i[31] la_oenb[0] wbs_adr_i[20] wbs_adr_i[21]
+ wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27]
+ wbs_adr_i[28] wbs_adr_i[29] la_oenb[1] wbs_adr_i[30] wbs_adr_i[31] la_oenb[2] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] la_oenb[3] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] la_oenb[4] wbs_dat_o[30] wbs_dat_o[31] la_oenb[5] la_data_in[0] la_data_in[1]
+ la_data_in[2] la_data_in[3] la_data_in[4] la_data_in[5] la_data_out[0] la_data_out[1]
+ la_data_out[2] la_data_out[3] la_data_out[4] la_data_out[5] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] la_data_in[26] la_data_in[11]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[6] la_data_in[7] la_data_in[8]
+ la_data_in[9] la_data_in[15] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_in[16] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[10]
+ la_data_out[6] la_data_out[7] la_data_out[8] la_data_out[9] la_data_in[20] la_oenb[10]
+ la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_data_in[21] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_data_in[22] la_data_in[39] la_oenb[45] la_data_in[40]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_in[41] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_in[42] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_oenb[46]
+ la_oenb[38] la_oenb[39] la_oenb[37] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_oenb[44] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_data_in[38] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[47] la_oenb[48]
+ la_oenb[49] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[60] la_data_in[61]
+ la_data_in[62] la_data_in[63] la_data_out[47] la_data_out[48] la_data_out[49] la_data_in[64]
+ la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_in[65] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_in[66] la_data_in[67] la_data_in[72]
+ la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78]
+ la_data_in[79] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[69] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_data_out[68] la_data_out[69]
+ la_data_in[70] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_in[71] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_in[68] la_oenb[88] la_oenb[89]
+ la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96]
+ la_oenb[97] la_oenb[98] la_oenb[99] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[100] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94]
+ la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[93] la_data_out[106] la_data_out[94] la_data_out[107] la_data_out[95]
+ la_data_out[96] la_data_out[108] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[92] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_data_in[88] la_data_in[89] la_data_out[88]
+ la_data_out[89] la_data_out[90] la_data_out[91] la_data_in[119] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_in[116] la_data_in[117] la_data_out[123]
+ la_data_in[112] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_in[118] la_oenb[109] la_data_in[120] la_oenb[110] la_data_in[121] la_oenb[111]
+ la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118]
+ la_oenb[119] la_data_in[122] la_data_in[123] la_oenb[120] la_oenb[121] la_oenb[122]
+ la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_out[110] user_clock2 user_irq[0]
+ la_data_in[113] user_irq[1] la_data_in[114] user_irq[2] la_data_out[111] la_data_out[112]
+ la_data_out[109] la_data_in[109] la_data_out[113] la_data_in[110] la_data_out[114]
+ la_oenb[108] la_data_out[115] la_data_out[116] la_data_in[111] la_data_out[117]
+ la_data_in[115] la_data_out[118] la_data_out[119] io_analog[4] io_analog[5] io_analog[6]
+ gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5] gpio_analog[6] gpio_noesd[2]
+ gpio_noesd[3] gpio_noesd[4] gpio_noesd[5] gpio_noesd[6] io_analog[0] io_analog[1]
+ io_analog[2] io_analog[3] io_clamp_high[0] io_clamp_low[0] io_in[10] io_in[11] io_in[12]
+ io_in[13] io_in[9] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12] io_in_3v3[13] io_in_3v3[9]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[9] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[9] vccd1 vdda1 vssa1 io_in[16] io_in[17] gpio_analog[9] gpio_noesd[10]
+ io_analog[7] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_analog[8]
+ io_analog[9] gpio_noesd[7] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] gpio_noesd[8]
+ io_clamp_high[1] io_clamp_high[2] gpio_noesd[9] io_clamp_low[1] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_clamp_low[2] gpio_analog[10] io_analog[10] vccd2 gpio_analog[7]
+ gpio_analog[8] io_in[14] io_in[15] vssa2 io_in_3v3[24] io_in_3v3[25] io_in_3v3[26]
+ gpio_analog[16] gpio_analog[17] gpio_analog[11] gpio_analog[12] gpio_noesd[11] io_in[18]
+ io_in[19] io_in[20] io_in[21] io_oeb[18] io_oeb[19] io_oeb[20] io_oeb[21] io_oeb[22]
+ io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] io_out[18]
+ io_out[19] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26]
+ gpio_noesd[16] gpio_noesd[17] gpio_analog[13] gpio_analog[14] gpio_analog[15] io_in_3v3[18]
+ io_in_3v3[19] vdda2 io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23] vssd2
+ io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in[1] io_oeb[0] gpio_noesd[0] io_in[2]
+ io_in[3] io_in[4] io_in[5] io_out[1] io_in[6] io_in_3v3[1] io_in[7] io_in[8] gpio_analog[0]
+ io_oeb[1] io_in_3v3[0] io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] gpio_analog[1] gpio_noesd[1] io_in[0] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] vssd1 io_in_3v3[5]
+ io_out[0]
Xesd_diodes_0 vccd2 io_analog[10] vssd2 dw_10605_683750# esd_diodes
Xesd_diodes_1 vccd2 io_analog[9] vssd2 dw_10605_686997# esd_diodes
XVGA_final_0 io_analog[8] io_analog[7] VGA_final_0/RF_in VGA_final_0/RF_out io_analog[5]
+ io_analog[6] VGA_final
Xesd_0 vdda1 io_analog[0] dw_514926_556356# dw_510516_556356# esd_0/out vssa1 esd
XCascode_Amp_0 Cascode_Amp_0/Vgg_1v8 Cascode_Amp_0/RF_out Cascode_Amp_0/RF_in Cascode_Amp_0/gnd
+ Cascode_Amp
XCascode_Amp_1 Cascode_Amp_1/Vgg_1v8 Cascode_Amp_1/RF_out Cascode_Amp_1/RF_in Cascode_Amp_1/gnd
+ Cascode_Amp
Xsar_adc_0 io_analog[9] io_analog[10] io_out[24] io_in[25] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[20] io_out[21] io_out[22] io_out[23] io_in[26]
+ vccd2 vssd2 sar_adc
XLNA_final_0 io_analog[3] LNA_final_0/RF_in LNA_final_0/RF_out io_analog[2] io_analog[4]
+ LNA_final
Xfull_IC_1_0 esd_0/out out_buf_0/in vdda1 io_in[8] io_in[9] io_in[10] io_in[11] io_in[12]
+ io_out[13] vssa1 full_IC_1
XStandalone_mosfet_32f_0 Standalone_mosfet_32f_0/signal_out Standalone_mosfet_32f_0/signal_in
+ Standalone_mosfet_32f_0/gnd Standalone_mosfet_32f
XStandalone_mosfet_32f_1 Standalone_mosfet_32f_1/signal_out Standalone_mosfet_32f_1/signal_in
+ Standalone_mosfet_32f_1/gnd Standalone_mosfet_32f
XRF_switch_0 gpio_analog[0] RF_switch_0/Port3 RF_switch_0/Port1 RF_switch_0/Port2
+ vdda1 vssd1 RF_switch
Xout_buf_0 out_buf_0/in io_analog[1] vdda1 vssa1 out_buf
XStandalone_mosfet_150f_0 Standalone_mosfet_150f_0/signal_in Standalone_mosfet_150f_0/signal_out
+ Standalone_mosfet_150f_0/gnd Standalone_mosfet_150f
XStandalone_mosfet_150f_1 Standalone_mosfet_150f_1/signal_in Standalone_mosfet_150f_1/signal_out
+ Standalone_mosfet_150f_1/gnd Standalone_mosfet_150f
R0 vssa1 vssd1 sky130_fd_pr__res_generic_m3 w=3.635e+07u l=1.7e+07u
.ends

